../ip_repo/accelerator_1.0/src/user_app.vhd