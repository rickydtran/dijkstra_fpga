../ip_repo/accelerator_1.0/src/config_pkg.vhd