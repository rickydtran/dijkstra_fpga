../ip_repo/accelerator_1.0/src/add_pipe.vhd