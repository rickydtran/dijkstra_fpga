../ip_repo/accelerator_1.0/src/memory_map.vhd