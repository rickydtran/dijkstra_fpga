../ip_repo/accelerator_1.0/src/ctrl.vhd