-- Ricky Tran
-- University of Florida
-- user_app_tb.vhd

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.config_pkg.all;
use work.user_pkg.all;

entity user_app_tb is
end user_app_tb;

architecture tb of user_app_tb is
  type t_2d_a is array(0 to 63, 0 to 63) of integer range 0 to 255;
  constant input_key : t_2d_a :=
  ((    0,   238,    35,   209,   219,    61,    35,    94,     7,   251,   157,   245,    42,   114,   117,    33,     8,   102,   153,   187,     7,     1,    47,   185,    43,    63,    14,    84,    31,   246,   127,   249,    35,   119,    65,     0,   233,   109,     0,   218,   166,    56,   145,    22,    45,   129,    80,    26,   180,    77,   214,   160,    28,     0,    13,   165,     0,   114,   191,    50,    88,   142,    44,     8),
   (  238,     0,   234,    26,    10,    63,     0,   225,   109,   197,   212,   184,    57,   255,    56,    54,   237,     0,    47,     0,   207,   154,   154,   103,     7,     0,   240,   226,    13,   180,    19,   124,    61,   251,   154,   211,    60,    74,     8,     0,    24,   219,   253,   227,    32,   167,   142,     0,   121,   178,   180,   239,    24,     0,   161,   184,   167,    91,     2,     0,    12,    19,     0,    24),
   (   35,   234,     0,     0,   238,   128,   190,     0,   160,   137,   185,   131,   228,    56,    59,   211,    12,    67,   212,     5,    13,   186,    80,   236,   190,   209,     0,   191,     0,   252,   248,    90,    12,   102,    44,   195,    20,    42,     0,   201,     5,    27,     0,     6,     0,    15,    89,   142,    27,    59,    28,   219,   198,    16,   211,    89,    16,   128,   245,    87,   130,    83,   128,     0),
   (  209,    26,     0,     0,   188,   142,     0,     8,   169,   114,   153,   206,   138,   105,    19,    78,    72,    30,   224,    93,    67,    69,   229,   139,   122,    31,    90,   144,    14,     0,    25,   150,    15,   208,     0,    37,   180,    39,   110,   247,    16,   211,    24,    69,    15,    54,    40,   219,     0,   206,   208,    40,   140,   167,    97,     0,     6,   246,   182,   221,   185,     0,   126,     0),
   (  219,    10,   238,   188,     0,    20,    42,   196,    32,   120,    30,   233,   210,    55,   100,   245,   172,   170,    52,   194,   170,   129,    42,    92,   145,     0,   226,   219,   238,    57,   194,   226,    22,   173,   127,   116,   110,    70,     0,   155,   141,    95,   239,    15,    21,   155,   191,    82,    13,    48,     0,    20,   165,    42,   146,    30,   139,    37,   156,    99,   220,    47,    59,   188),
   (   61,    63,   128,   142,    20,     0,   132,   205,   156,   154,    60,     0,    94,   254,   108,    37,   196,   249,    42,   102,   179,   141,   213,   214,   240,    33,   115,    58,    66,   235,   108,   169,    49,   224,   232,   151,   160,   131,     0,   197,   172,     0,   200,   253,   154,    20,    83,   126,     0,   236,   109,   235,   137,   242,   211,     0,    95,   148,   179,   225,    86,    13,    14,    13),
   (   35,     0,   190,     0,    42,   132,     0,   150,    12,   202,     0,   148,   230,   163,   124,   167,   213,    71,    44,   103,    63,    11,    78,     0,   162,   122,   224,   159,   223,   208,   177,   182,   249,    23,   241,    73,   112,   225,   141,   169,     5,   198,   145,   188,     0,    94,   127,   173,   224,   124,   163,    30,    46,    14,   155,   164,   120,    89,   222,    69,   106,   211,   212,     0),
   (   94,   225,     0,     8,   196,   205,   150,     0,   183,    22,    78,    67,   206,    56,   105,   137,    34,   163,   199,   178,    10,   223,   250,    82,    16,   199,   138,    33,   110,    62,    69,   199,    98,   113,    68,    15,    74,   143,   245,   194,    15,    93,   187,   229,    58,   165,    53,     5,   138,   229,   226,   117,    36,     0,   178,     0,   210,   198,    94,   221,    83,   175,    33,   233),
   (    7,   109,   160,   169,    32,   156,    12,   183,     0,   156,   223,   178,   208,   127,    35,   162,   126,    89,   138,   196,   236,    33,   151,    90,    64,    36,    18,   107,   150,    48,   255,   242,   141,    67,    25,   194,   184,    93,   101,   121,   247,    65,   144,   201,   173,   135,    11,    71,   225,   184,   107,   244,    50,   168,   205,     0,   241,    67,    25,   139,     0,   198,   180,   248),
   (  251,   197,   137,   114,   120,   154,   202,    22,   156,     0,   158,   203,    76,    40,    90,    77,    59,    86,    54,   133,   116,   136,     0,     0,   186,    65,   241,    53,   177,   185,     0,    67,   238,   243,    48,   214,   212,   145,     7,   250,   250,     6,     0,     8,    26,   171,   218,    43,    26,   232,   131,    50,   206,   213,    92,   241,   134,     0,   208,    83,    56,    14,   163,   156),
   (  157,   212,   185,   153,    30,    60,     0,    78,   223,   158,     0,   143,    65,   159,   241,   134,    14,   215,    61,   150,   238,   232,    41,    19,   201,   142,   210,    71,   158,     1,    62,    58,     0,   208,   225,     0,   175,    90,     4,     0,   201,   233,   197,    34,    97,   167,   146,     0,    60,    81,    55,   225,    69,   239,   111,    93,    74,     0,    91,   254,   192,   147,   178,   191),
   (  245,   184,   131,   206,   233,     0,   148,    67,   178,   203,   143,     0,    87,    89,    71,     0,    81,    32,     0,   249,    63,   201,   203,   216,   178,    97,   234,   118,   131,   145,    71,   137,   247,     0,   111,     0,   214,     0,    93,   243,   177,    99,   215,    27,    35,    98,   100,    96,   191,    96,    56,    49,   222,    69,   129,   137,   131,   174,   159,    99,    19,   137,    52,     0),
   (   42,    57,   228,   138,   210,    94,   230,   206,   208,    76,    65,    87,     0,   178,   247,   215,   238,     0,    60,   180,    89,    19,   150,   242,    69,    21,   165,    66,    83,   207,    14,    77,   199,   168,   246,   160,    91,   197,   150,   106,     0,   201,    87,   128,   114,   226,    27,   154,   157,   136,    76,   207,    96,   163,    86,    48,   196,   211,     0,   186,   230,   182,   248,    72),
   (  114,   255,    56,   105,    55,   254,   163,    56,   127,    40,   159,    89,   178,     0,    66,   232,   133,     7,    14,   117,   216,    40,   165,     9,   243,   182,    85,   214,   164,   168,    72,   106,    42,    46,    17,   155,     8,    20,   161,   195,   115,    36,     0,    21,   230,   129,   241,     0,    96,    61,    90,    73,   118,   253,   171,     0,    54,   222,   219,   244,   109,     0,    57,   137),
   (  117,    56,    59,    19,   100,   108,   124,   105,    35,    90,   241,    71,   247,    66,     0,   218,   155,   206,    42,   183,   214,   178,   102,    46,    49,   250,   145,   119,    64,   172,     0,   134,   237,   142,   213,   249,     0,    25,   238,    97,     8,    12,   248,    17,    58,   194,    29,   155,   169,    19,     8,   224,    85,   254,   184,   243,    92,   126,    87,    84,   144,    25,   155,   144),
   (   33,    54,   211,    78,   245,    37,   167,   137,   162,    77,   134,     0,   215,   232,   218,     0,    17,   118,     0,   144,   164,    23,    91,   171,    23,   113,     0,     0,   211,   151,    64,   151,    59,   191,   108,    75,   211,     0,   119,     2,   116,     0,    38,   204,   212,    52,   241,   163,    18,   219,   238,   199,   101,     0,    28,    40,   203,     0,   141,    29,   197,   184,   140,     0),
   (    8,   237,    12,    72,   172,   196,   213,    34,   126,    59,    14,    81,   238,   133,   155,    17,     0,    12,   158,    52,    56,     0,   249,   112,    26,   187,    82,   228,    99,    19,   198,   201,   118,   209,    30,   212,   194,   122,   243,   237,    23,   115,    78,   116,   230,    54,    26,    94,    90,     0,   135,   183,   210,   135,   126,    81,   240,     0,   168,   144,   146,   164,   182,   230),
   (  102,     0,    67,    30,   170,   249,    71,   163,    89,    86,   215,    32,     0,     7,   206,   118,    12,     0,     0,     4,     0,   192,   215,   174,     0,   148,   216,   208,    80,     0,   233,    58,    64,   122,   199,   169,   246,   228,   121,     0,   178,    79,   142,   166,   166,    59,   226,   136,    10,   206,    64,   203,    97,   139,    49,    87,   148,     8,   113,    67,    93,    93,    30,    32),
   (  153,    47,   212,   224,    52,    42,    44,   199,   138,    54,    61,     0,    60,    14,    42,     0,   158,     0,     0,    45,   195,   237,    24,     0,    72,   208,   108,     0,    46,   147,    90,    45,   183,    61,   128,    71,   127,   233,   146,   130,    18,    64,    59,   235,     0,   204,   207,    46,   231,   254,     0,    84,   229,    70,   238,    35,   111,    84,   235,    97,   205,   117,   128,   144),
   (  187,     0,     5,    93,   194,   102,   103,   178,   196,   133,   150,   249,   180,   117,   183,   144,    52,     4,    45,     0,    31,     0,    15,   102,     0,   228,   210,    28,     0,   118,   203,   226,    84,    19,   180,   242,   161,    50,   230,    59,   173,    39,   116,    58,    93,    17,   112,    20,   203,   168,   221,    72,     0,    20,   157,   121,   205,   168,   103,   102,    53,    87,    53,    16),
   (    7,   207,    13,    67,   170,   179,    63,    10,   236,   116,   238,    63,    89,   216,   214,   164,    56,     0,   195,    31,     0,    80,   192,    27,   178,    52,   150,    49,     0,     0,   185,   102,   225,   180,   144,     0,   108,   203,   244,   240,   137,     0,   144,    88,     0,     4,   161,   193,   212,    63,   184,   179,   246,   167,    71,   224,   164,   127,   172,    74,    17,   216,   214,   173),
   (    1,   154,   186,    69,   129,   141,    11,   223,    33,   136,   232,   201,    19,    40,   178,    23,     0,   192,   237,     0,    80,     0,    10,    85,    45,    24,   249,    95,   163,   147,   224,    13,    42,   205,    26,     8,    91,   124,   148,    74,     0,    69,     0,    80,    63,     0,    92,   233,   166,   135,   169,    76,    72,   237,   173,    22,   147,    18,    31,   195,   178,    75,   124,   119),
   (   47,   154,    80,   229,    42,   213,    78,   250,   151,     0,    41,   203,   150,   165,   102,    91,   249,   215,    24,    15,   192,    10,     0,    31,   204,   172,   149,   160,   140,    79,     0,    66,   143,    27,     0,   207,     0,     0,    16,   230,   190,    76,   133,   143,    32,   205,   208,   176,   205,   136,   118,   147,   227,   201,   161,   154,   234,    99,    79,   100,    93,    93,   141,    23),
   (  185,   103,   236,   139,    92,   214,     0,    82,    90,     0,    19,   216,   242,     9,    46,   171,   112,   174,     0,   102,    27,    85,    31,     0,    29,   238,   193,     0,    22,   133,    38,    74,    32,    48,   224,   165,     0,   236,   183,   253,   158,   207,     0,   235,   188,   229,     0,   249,   204,    47,     0,    53,    47,     9,   118,    71,   237,   132,    41,   111,    94,    41,   166,    57),
   (   43,     7,   190,   122,   145,   240,   162,    16,    64,   186,   201,   178,    69,   243,    49,    23,    26,     0,    72,     0,   178,    45,   204,    29,     0,    57,     0,   222,    35,    37,   247,   190,    20,   204,   217,     2,   177,    12,   213,   194,   136,    66,    48,   133,     0,     0,    92,   246,    16,   133,   205,    84,    46,   169,   112,     6,   232,    89,    31,   146,    60,   242,    55,   222),
   (   63,     0,   209,    31,     0,    33,   122,   199,    36,    65,   142,    97,    21,   182,   250,   113,   187,   148,   208,   228,    52,    24,   172,   238,    57,     0,   166,   220,   225,     0,   105,   209,   128,    44,    19,    32,   132,   227,   199,     0,   138,    50,    49,    88,     6,   101,    84,   218,   182,    17,   255,     0,    48,    88,   159,     0,     2,   144,   171,    74,   202,    17,    11,     0),
   (   14,   240,     0,    90,   226,   115,   224,   138,    18,   241,   210,   234,   165,    85,   145,     0,    82,   216,   108,   210,   150,   249,   149,   193,     0,   166,     0,   250,   202,   110,   146,   167,   231,     9,   123,   145,    64,     0,   238,    55,    31,   136,    89,   222,   123,   106,    68,   220,    87,    82,   233,   209,   169,    22,     3,     0,    36,     4,    24,    92,    97,    84,   184,    45),
   (   84,   226,   191,   144,   219,    58,   159,    33,   107,    53,    71,   118,    66,   214,   119,     0,   228,   208,     0,    28,    49,    95,   160,     0,   222,   220,   250,     0,    39,   121,     0,    37,   200,   133,    49,   112,   150,     0,   114,   227,   230,   156,   104,   129,    21,   104,   139,   111,    24,   110,   122,    63,   245,   110,   168,     0,     5,    10,    84,   198,   216,     0,   145,   148),
   (   31,    13,     0,    14,   238,    66,   223,   110,   150,   177,   158,   131,    83,   164,    64,   211,    99,    80,    46,     0,     0,   163,   140,    22,    35,   225,   202,    39,     0,     0,    44,   140,   170,   149,   226,    26,    36,   204,    43,    20,    30,    14,   234,    55,   163,   123,   187,    51,   151,    19,    28,   110,    91,    50,    40,   236,     0,    72,    70,   109,   226,   126,   197,    99),
   (  246,   180,   252,     0,    57,   235,   208,    62,    48,   185,     1,   145,   207,   168,   172,   151,    19,     0,   147,   118,     0,   147,    79,   133,    37,     0,   110,   121,     0,     0,    23,    86,    56,   209,    71,   105,   252,   202,   127,   132,    64,    73,    26,    46,   236,   154,     8,   131,    47,   224,    43,    59,    54,     0,   225,   159,    42,   102,     9,   183,    56,     5,     3,   116),
   (  127,    19,   248,    25,   194,   108,   177,    69,   255,     0,    62,    71,    14,    72,     0,    64,   198,   233,    90,   203,   185,   224,     0,    38,   247,   105,   146,     0,    44,    23,     0,   121,   188,    21,   155,   248,   180,   212,   118,    25,    14,   100,    66,    97,   141,    56,   108,     0,   168,   240,   155,    15,    66,   212,     0,   195,    16,    36,   190,   254,   181,     0,    78,     0),
   (  249,   124,    90,   150,   226,   169,   182,   199,   242,    67,    58,   137,    77,   106,   134,   151,   201,    58,    45,   226,   102,    13,    66,    74,   190,   209,   167,    37,   140,    86,   121,     0,     9,   156,   159,   172,   195,   224,    52,    65,   225,    20,    83,   137,   126,    18,   243,   233,   146,   145,   226,   104,    72,   206,   140,   124,    38,   127,   203,    71,   133,   126,   122,    65),
   (   35,    61,    12,    15,    22,    49,   249,    98,   141,   238,     0,   247,   199,    42,   237,    59,   118,    64,   183,    84,   225,    42,   143,    32,    20,   128,   231,   200,   170,    56,   188,     9,     0,    89,   107,   135,   109,   201,     0,    95,   111,    65,     7,   186,   127,   121,   234,   211,    61,    30,   102,    35,    46,    58,   215,    70,     0,    24,   155,   113,   130,    56,   221,   201),
   (  119,   251,   102,   208,   173,   224,    23,   113,    67,   243,   208,     0,   168,    46,   142,   191,   209,   122,    61,    19,   180,   205,    27,    48,   204,    44,     9,   133,   149,   209,    21,   156,    89,     0,   124,   153,   135,   249,   226,   162,   140,     0,    62,   162,   173,   154,     0,   191,   198,   207,    97,     0,   214,    32,    95,    42,   175,   141,   106,    15,   204,    86,   203,   233),
   (   65,   154,    44,     0,   127,   232,   241,    68,    25,    48,   225,   111,   246,    17,   213,   108,    30,   199,   128,   180,   144,    26,     0,   224,   217,    19,   123,    49,   226,    71,   155,   159,   107,   124,     0,   100,    76,    57,   185,     3,    17,    91,    59,   208,    60,    88,    51,     8,     0,    14,   196,   153,   126,    56,    21,     0,   186,   157,   206,   195,   254,   176,   117,    17),
   (    0,   211,   195,    37,   116,   151,    73,    15,   194,   214,     0,     0,   160,   155,   249,    75,   212,   169,    71,   242,     0,     8,   207,   165,     2,    32,   145,   112,    26,   105,   248,   172,   135,   153,   100,     0,    54,   197,   181,   255,   238,   218,   251,   235,   106,    35,   180,    89,   215,   205,   106,   115,   146,   226,    29,    33,     4,   159,   231,    82,    58,   191,   192,   215),
   (  233,    60,    20,   180,   110,   160,   112,    74,   184,   212,   175,   214,    91,     8,     0,   211,   194,   246,   127,   161,   108,    91,     0,     0,   177,   132,    64,   150,    36,   252,   180,   195,   109,   135,    76,    54,     0,     4,    96,    15,     8,    29,    80,   115,   213,     0,    23,    84,   221,    79,   243,   201,   189,   234,   119,    59,    33,    54,   220,   125,   187,    87,   204,   209),
   (  109,    74,    42,    39,    70,   131,   225,   143,    93,   145,    90,     0,   197,    20,    25,     0,   122,   228,   233,    50,   203,   124,     0,   236,    12,   227,     0,     0,   204,   202,   212,   224,   201,   249,    57,   197,     4,     0,   209,    50,    13,    80,    99,   246,   172,    50,   136,   218,    47,   248,   160,   223,   169,    70,   134,   187,   239,   255,    34,   158,     0,   152,   182,   190),
   (    0,     8,     0,   110,     0,     0,   141,   245,   101,     7,     4,    93,   150,   161,   238,   119,   243,   121,   146,   230,   244,   148,    16,   183,   213,   199,   238,   114,    43,   127,   118,    52,     0,   226,   185,   181,    96,   209,     0,     0,    46,    91,   149,    83,   100,   168,     1,   180,   112,    56,     0,   144,   129,   243,   117,   232,    50,   150,    30,   220,    10,   180,   233,   103),
   (  218,     0,   201,   247,   155,   197,   169,   194,   121,   250,     0,   243,   106,   195,    97,     2,   237,     0,   130,    59,   240,    74,   230,   253,   194,     0,    55,   227,    20,   132,    25,    65,    95,   162,     3,   255,    15,    50,     0,     0,   150,   231,   131,    21,   227,   168,    23,   166,   180,    69,     0,     0,   124,   254,   152,    57,   232,   235,   167,    38,     0,    31,    75,    55),
   (  166,    24,     5,    16,   141,   172,     5,    15,   247,   250,   201,   177,     0,   115,     8,   116,    23,   178,    18,   173,   137,     0,   190,   158,   136,   138,    31,   230,    30,    64,    14,   225,   111,   140,    17,   238,     8,    13,    46,   150,     0,     0,    27,    71,     7,   236,   135,   231,     0,    44,    31,     0,   212,    87,   193,    83,    54,   239,     0,    47,     0,    77,   163,   122),
   (   56,   219,    27,   211,    95,     0,   198,    93,    65,     6,   233,    99,   201,    36,    12,     0,   115,    79,    64,    39,     0,    69,    76,   207,    66,    50,   136,   156,    14,    73,   100,    20,    65,     0,    91,   218,    29,    80,    91,   231,     0,     0,   141,     0,   178,    55,   204,   139,    12,   254,     0,   171,   128,    54,    79,   214,   160,     0,    78,     5,    17,   109,     0,   106),
   (  145,   253,     0,    24,   239,   200,   145,   187,   144,     0,   197,   215,    87,     0,   248,    38,    78,   142,    59,   116,   144,     0,   133,     0,    48,    49,    89,   104,   234,    26,    66,    83,     7,    62,    59,   251,    80,    99,   149,   131,    27,   141,     0,    56,    78,   154,   164,    10,   179,    93,    31,   174,    32,     0,    52,    43,   118,   147,   159,   154,     0,     4,     5,   218),
   (   22,   227,     6,    69,    15,   253,   188,   229,   201,     8,    34,    27,   128,    21,    17,   204,   116,   166,   235,    58,    88,    80,   143,   235,   133,    88,   222,   129,    55,    46,    97,   137,   186,   162,   208,   235,   115,   246,    83,    21,    71,     0,    56,     0,    44,    17,    67,    60,    11,     5,   119,   134,   132,   209,    89,   251,    40,   176,    42,   103,   143,    64,   228,   182),
   (   45,    32,     0,    15,    21,   154,     0,    58,   173,    26,    97,    35,   114,   230,    58,   212,   230,   166,     0,    93,     0,    63,    32,   188,     0,     6,   123,    21,   163,   236,   141,   126,   127,   173,    60,   106,   213,   172,   100,   227,     7,   178,    78,    44,     0,   192,   208,    49,     0,     0,   108,   193,   255,   253,    21,   128,   187,   241,     0,   193,    98,    39,   182,     1),
   (  129,   167,    15,    54,   155,    20,    94,   165,   135,   171,   167,    98,   226,   129,   194,    52,    54,    59,   204,    17,     4,     0,   205,   229,     0,   101,   106,   104,   123,   154,    56,    18,   121,   154,    88,    35,     0,    50,   168,   168,   236,    55,   154,    17,   192,     0,   249,   115,     0,    93,   132,    36,     0,   117,   148,    69,    90,     0,   127,   248,   244,   186,   153,   112),
   (   80,   142,    89,    40,   191,    83,   127,    53,    11,   218,   146,   100,    27,   241,    29,   241,    26,   226,   207,   112,   161,    92,   208,     0,    92,    84,    68,   139,   187,     8,   108,   243,   234,     0,    51,   180,    23,   136,     1,    23,   135,   204,   164,    67,   208,   249,     0,    26,   192,   138,    65,   108,    69,   180,    67,   155,    77,   125,    39,   124,   203,   237,    39,   126),
   (   26,     0,   142,   219,    82,   126,   173,     5,    71,    43,     0,    96,   154,     0,   155,   163,    94,   136,    46,    20,   193,   233,   176,   249,   246,   218,   220,   111,    51,   131,     0,   233,   211,   191,     8,    89,    84,   218,   180,   166,   231,   139,    10,    60,    49,   115,    26,     0,   166,    44,    45,   252,   203,   105,   170,    23,    89,   243,    90,    11,   111,   203,   224,   250),
   (  180,   121,    27,     0,    13,     0,   224,   138,   225,    26,    60,   191,   157,    96,   169,    18,    90,    10,   231,   203,   212,   166,   205,   204,    16,   182,    87,    24,   151,    47,   168,   146,    61,   198,     0,   215,   221,    47,   112,   180,     0,    12,   179,    11,     0,     0,   192,   166,     0,     0,     0,    73,    80,    49,    84,    89,    21,     0,   185,     4,   249,    99,     0,     0),
   (   77,   178,    59,   206,    48,   236,   124,   229,   184,   232,    81,    96,   136,    61,    19,   219,     0,   206,   254,   168,    63,   135,   136,    47,   133,    17,    82,   110,    19,   224,   240,   145,    30,   207,    14,   205,    79,   248,    56,    69,    44,   254,    93,     5,     0,    93,   138,    44,     0,     0,   180,     0,   194,   134,    53,    41,   161,   160,   214,   137,   180,    67,   176,   180),
   (  214,   180,    28,   208,     0,   109,   163,   226,   107,   131,    55,    56,    76,    90,     8,   238,   135,    64,     0,   221,   184,   169,   118,     0,   205,   255,   233,   122,    28,    43,   155,   226,   102,    97,   196,   106,   243,   160,     0,     0,    31,     0,    31,   119,   108,   132,    65,    45,     0,   180,     0,   229,   117,   179,   231,    25,     0,     0,     1,   107,   215,   113,    56,   226),
   (  160,   239,   219,    40,    20,   235,    30,   117,   244,    50,   225,    49,   207,    73,   224,   199,   183,   203,    84,    72,   179,    76,   147,    53,    84,     0,   209,    63,   110,    59,    15,   104,    35,     0,   153,   115,   201,   223,   144,     0,     0,   171,   174,   134,   193,    36,   108,   252,    73,     0,   229,     0,   109,   225,    81,   106,   221,   242,   238,   192,   246,    26,    26,   194),
   (   28,    24,   198,   140,   165,   137,    46,    36,    50,   206,    69,   222,    96,   118,    85,   101,   210,    97,   229,     0,   246,    72,   227,    47,    46,    48,   169,   245,    91,    54,    66,    72,    46,   214,   126,   146,   189,   169,   129,   124,   212,   128,    32,   132,   255,     0,    69,   203,    80,   194,   117,   109,     0,   142,   116,   136,   153,    27,   178,   196,     0,   204,    84,    93),
   (    0,     0,    16,   167,    42,   242,    14,     0,   168,   213,   239,    69,   163,   253,   254,     0,   135,   139,    70,    20,   167,   237,   201,     9,   169,    88,    22,   110,    50,     0,   212,   206,    58,    32,    56,   226,   234,    70,   243,   254,    87,    54,     0,   209,   253,   117,   180,   105,    49,   134,   179,   225,   142,     0,   164,   246,   131,    66,   130,   119,   187,   247,    43,    45),
   (   13,   161,   211,    97,   146,   211,   155,   178,   205,    92,   111,   129,    86,   171,   184,    28,   126,    49,   238,   157,    71,   173,   161,   118,   112,   159,     3,   168,    40,   225,     0,   140,   215,    95,    21,    29,   119,   134,   117,   152,   193,    79,    52,    89,    21,   148,    67,   170,    84,    53,   231,    81,   116,   164,     0,    20,    87,    78,   156,    95,     4,     0,   196,    44),
   (  165,   184,    89,     0,    30,     0,   164,     0,     0,   241,    93,   137,    48,     0,   243,    40,    81,    87,    35,   121,   224,    22,   154,    71,     6,     0,     0,     0,   236,   159,   195,   124,    70,    42,     0,    33,    59,   187,   232,    57,    83,   214,    43,   251,   128,    69,   155,    23,    89,    41,    25,   106,   136,   246,    20,     0,    47,    95,    45,   145,   226,    64,    92,   247),
   (    0,   167,    16,     6,   139,    95,   120,   210,   241,   134,    74,   131,   196,    54,    92,   203,   240,   148,   111,   205,   164,   147,   234,   237,   232,     2,    36,     5,     0,    42,    16,    38,     0,   175,   186,     4,    33,   239,    50,   232,    54,   160,   118,    40,   187,    90,    77,    89,    21,   161,     0,   221,   153,   131,    87,    47,     0,   195,   147,    69,   159,   113,   249,    67),
   (  114,    91,   128,   246,    37,   148,    89,   198,    67,     0,     0,   174,   211,   222,   126,     0,     0,     8,    84,   168,   127,    18,    99,   132,    89,   144,     4,    10,    72,   102,    36,   127,    24,   141,   157,   159,    54,   255,   150,   235,   239,     0,   147,   176,   241,     0,   125,   243,     0,   160,     0,   242,    27,    66,    78,    95,   195,     0,   144,    66,   226,    39,    88,    28),
   (  191,     2,   245,   182,   156,   179,   222,    94,    25,   208,    91,   159,     0,   219,    87,   141,   168,   113,   235,   103,   172,    31,    79,    41,    31,   171,    24,    84,    70,     9,   190,   203,   155,   106,   206,   231,   220,    34,    30,   167,     0,    78,   159,    42,     0,   127,    39,    90,   185,   214,     1,   238,   178,   130,   156,    45,   147,   144,     0,    21,    26,   126,   157,    30),
   (   50,     0,    87,   221,    99,   225,    69,   221,   139,    83,   254,    99,   186,   244,    84,    29,   144,    67,    97,   102,    74,   195,   100,   111,   146,    74,    92,   198,   109,   183,   254,    71,   113,    15,   195,    82,   125,   158,   220,    38,    47,     5,   154,   103,   193,   248,   124,    11,     4,   137,   107,   192,   196,   119,    95,   145,    69,    66,    21,     0,    28,   121,    89,     8),
   (   88,    12,   130,   185,   220,    86,   106,    83,     0,    56,   192,    19,   230,   109,   144,   197,   146,    93,   205,    53,    17,   178,    93,    94,    60,   202,    97,   216,   226,    56,   181,   133,   130,   204,   254,    58,   187,     0,    10,     0,     0,    17,     0,   143,    98,   244,   203,   111,   249,   180,   215,   246,     0,   187,     4,   226,   159,   226,    26,    28,     0,   118,     0,    22),
   (  142,    19,    83,     0,    47,    13,   211,   175,   198,    14,   147,   137,   182,     0,    25,   184,   164,    93,   117,    87,   216,    75,    93,    41,   242,    17,    84,     0,   126,     5,     0,   126,    56,    86,   176,   191,    87,   152,   180,    31,    77,   109,     4,    64,    39,   186,   237,   203,    99,    67,   113,    26,   204,   247,     0,    64,   113,    39,   126,   121,   118,     0,   196,   165),
   (   44,     0,   128,   126,    59,    14,   212,    33,   180,   163,   178,    52,   248,    57,   155,   140,   182,    30,   128,    53,   214,   124,   141,   166,    55,    11,   184,   145,   197,     3,    78,   122,   221,   203,   117,   192,   204,   182,   233,    75,   163,     0,     5,   228,   182,   153,    39,   224,     0,   176,    56,    26,    84,    43,   196,    92,   249,    88,   157,    89,     0,   196,     0,   139),
   (    8,    24,     0,     0,   188,    13,     0,   233,   248,   156,   191,     0,    72,   137,   144,     0,   230,    32,   144,    16,   173,   119,    23,    57,   222,     0,    45,   148,    99,   116,     0,    65,   201,   233,    17,   215,   209,   190,   103,    55,   122,   106,   218,   182,     1,   112,   126,   250,     0,   180,   226,   194,    93,    45,    44,   247,    67,    28,    30,     8,    22,   165,   139,     0));
   
  type list is array(0 to 1842) of integer;
  constant edge_list : list :=
  ( 494, 1243, 1341, 1571, 2055, 2555, 2717, 3061, 3873, 4454, 4761, 5051, 5377, 5679, 6187, 6670, 6996, 8227, 8567, 9449, 11030, 12468, 13014, 13837, 14706, 15448, 15916, 16136, 17178, 17418, 18401, 19384, 19513, 20024, 20717, 22170, 22535, 23280, 23522, 23565, 24444, 24637, 25083, 25555, 25660, 26648, 27619, 27680, 28302, 28793, 29106, 29720, 30369, 31234, 32019, 32536, 32803, 33258, 34030, 34176, 34494, 34976, 35209, 35513, 35715, 36152, 36819, 37588, 38330, 39377, 40696, 40794, 40972, 42004, 42282, 42953, 43013, 45371, 46043, 47120, 47488, 48768, 49361, 50364, 51570, 51865, 52174, 52362, 52755, 53070, 53320, 53984, 54109, 54339, 54597, 55013, 55179, 55583, 55898, 56334, 57808, 58548, 58990, 59859, 60431, 62160, 63494, 63990, 64182, 64697, 67114, 67960, 68126, 68585, 68919, 69220, 69621, 69804, 70058, 70826, 71210, 71516, 73410, 74157, 74367, 74612, 74862, 75917, 76527, 76559, 77503, 77650, 77837, 78612, 79013, 79146, 79506, 81467, 81852, 82239, 82830, 82964, 84378, 84540, 85086, 85502, 85797, 86521, 86886, 87765, 88304, 88353, 90025, 90592, 90856, 91031, 91296, 91523, 92101, 92872, 93181, 94700, 95211, 95369, 95955, 96660, 97249, 97366, 97549, 97806, 98061, 99716, 100246, 100810, 101268, 102012, 102613, 103271, 103487, 103691, 104610, 105184, 105375, 105936, 106745, 107249, 107337, 107632, 108457, 108549, 108998, 109201, 109500, 109918, 110207, 110816, 111267, 112283, 112548, 113477, 114131, 114782, 115464, 115908, 116173, 116919, 117326, 117966, 118072, 119203, 119730, 120570, 121287, 121482, 121633, 122437, 122823, 122978, 123663, 123978, 124866, 124943, 125277, 126010, 126517, 127461, 127714, 127861, 128036, 129234, 129478, 130131, 130479, 130593, 131437, 132009, 132128, 132508, 132620, 134352, 134691, 135294, 135513, 136428, 136481, 137050, 137280, 137746, 138544, 139007, 139250, 139405, 140472, 140901, 141177, 141633, 141968, 142509, 144372, 144434, 144808, 145101, 145945, 146315, 147124, 147448, 147909, 149270, 149660, 150475, 151130, 151373, 151611, 151894, 152118, 152692, 154353, 154801, 155459, 155886, 156147, 157191, 157946, 157958, 158472, 158746, 159450, 159531, 159770, 160232, 160387, 160562, 161237, 162872, 163740, 164308, 166111, 166302, 166799, 167665, 167814, 168407, 168509, 168854, 169198, 169747, 170185, 170823, 171166, 171265, 171582, 173572, 174281, 174569, 174789, 174882, 175201, 175762, 176465, 177121, 177221, 177775, 179392, 179890, 182083, 182450, 183641, 184608, 186546, 187114, 187975, 189039, 191191, 191259, 191523, 192100, 192864, 193080, 193329, 193758, 194441, 194691, 195231, 195427, 196650, 197348, 197842, 198374, 198988, 199233, 199511, 200663, 201276, 201652, 201817, 202738, 203859, 204239, 205224, 205728, 205915, 207447, 207744, 208411, 209053, 209871, 210016, 210518, 210736, 211411, 211898, 212728, 213106, 213503, 213865, 214691, 215167, 215336, 215711, 216242, 217064, 217351, 217973, 218889, 219379, 219574, 219733, 220744, 221034, 221226, 221486, 222216, 222484, 222881, 223171, 223347, 223524, 224641, 226422, 226987, 227382, 227806, 228461, 228921, 229493, 229947, 230764, 231273, 232263, 232695, 232770, 233934, 234710, 235110, 235310, 235569, 236407, 236972, 237805, 238585, 238873, 239884, 240376, 240401, 241090, 241181, 241563, 242656, 242773, 243198, 243699, 243804, 244311, 244564, 245403, 246070, 247463, 247689, 247970, 249562, 251483, 251927, 253139, 253504, 254572, 254795, 255187, 255607, 255746, 256550, 256972, 257777, 258066, 258523, 259015, 259880, 260749, 260893, 261560, 261772, 262152, 262668, 263620, 263970, 264718, 265041, 265454, 265605, 265883, 266001, 266508, 267060, 267320, 268025, 268314, 269284, 269587, 270022, 270454, 270801, 271316, 271554, 272115, 272365, 272407, 272755, 272974, 273268, 274522, 275079, 275666, 275847, 276094, 276720, 277392, 277650, 278502, 279107, 279326, 280135, 282486, 283396, 286441, 286522, 286784, 287657, 287990, 288377, 289422, 289702, 290826, 291278, 291392, 291787, 293489, 293981, 294237, 295215, 295988, 296234, 296492, 296903, 297098, 298254, 298538, 299166, 299821, 300227, 300568, 301676, 302483, 302682, 302893, 303287, 304786, 305170, 305472, 305723, 306155, 306895, 306990, 307431, 308052, 308453, 308550, 308974, 309027, 309359, 309995, 310477, 311184, 311813, 312514, 313540, 313733, 314361, 315063, 315280, 318162, 318838, 319458, 320498, 321339, 321709, 322362, 322653, 322833, 323184, 323348, 324317, 325277, 325497, 326056, 326247, 326502, 327687, 328143, 328205, 329139, 329482, 330559, 331224, 331684, 332575, 333504, 333595, 334486, 335545, 336308, 336528, 337355, 338057, 338576, 338776, 339905, 340180, 340287, 340915, 341238, 341575, 341984, 342180, 342858, 343512, 343981, 344474, 345217, 345485, 346079, 346504, 346856, 347081, 347155, 347432, 347826, 347927, 348608, 348909, 349264, 350488, 350969, 351071, 351395, 351635, 351968, 352298, 352717, 352794, 353371, 353940, 355152, 356329, 356518, 356743, 357196, 358166, 359602, 361040, 362062, 362647, 363049, 363467, 363670, 363941, 365015, 365327, 365834, 366367, 366796, 367253, 367520, 367756, 367951, 368783, 368923, 369615, 370192, 370878, 371020, 371333, 371744, 372432, 372656, 373366, 373987, 374217, 374433, 375018, 375139, 376461, 376599, 377017, 377191, 377580, 378326, 378706, 379864, 380843, 381040, 381358, 381798, 382293, 383005, 383681, 384389, 385328, 385957, 386540, 386743, 387069, 387535, 388284, 388581, 389941, 390409, 390983, 391405, 391556, 392047, 392489, 392870, 393017, 393918, 394106, 394385, 395024, 395706, 396357, 397896, 398514, 398637, 399673, 400350, 400677, 401143, 401342, 402609, 403157, 404016, 404357, 405494, 405893, 406356, 406574, 407152, 407302, 407784, 408095, 408466, 408636, 409663, 411258, 411684, 411969, 412302, 412513, 412693, 413434, 413553, 413883, 414100, 414416, 414692, 414772, 415404, 415726, 416993, 417385, 417920, 418323, 418948, 419299, 419527, 419978, 420146, 420870, 421460, 422070, 422655, 422960, 423256, 423583, 423938, 424619, 425233, 427234, 427379, 428754, 429221, 429713, 430162, 430552, 432550, 433146, 433354, 433518, 434811, 435264, 436023, 436616, 436825, 437214, 437371, 437828, 438359, 438610, 439017, 439574, 440356, 440856, 441180, 441441, 442157, 443071, 443280, 443611, 443706, 444523, 444725, 445302, 445506, 445910, 446928, 447260, 447537, 448988, 450949, 452210, 452579, 452838, 453505, 453653, 453992, 454283, 454680, 455290, 455925, 456970, 457944, 458644, 458783, 460014, 460098, 460511, 460654, 460950, 461699, 462244, 462400, 462947, 463184, 463406, 464662, 464931, 465703, 466476, 466828, 467114, 468004, 469022, 469262, 469738, 469815, 470395, 470835, 471191, 471918, 472370, 472616, 473068, 473670, 473965, 474338, 474494, 474821, 475382, 475572, 475900, 476217, 476651, 476990, 477625, 478097, 478632, 479127, 482169, 482839, 483384, 484201, 484810, 485705, 486190, 486810, 486920, 487299, 487471, 488251, 489185, 489375, 489514, 489993, 490423, 490552, 490757, 491011, 491647, 491795, 492313, 492908, 493233, 494606, 496587, 497446, 498322, 499577, 499989, 500379, 500728, 501529, 502116, 502625, 502925, 503404, 504475, 504591, 504898, 505795, 505872, 506878, 507061, 507470, 508153, 508822, 509154, 509622, 510522, 510857, 511053, 511622, 511895, 512201, 513126, 513293, 513602, 513866, 514513, 514727, 514853, 515414, 516105, 516508, 516767, 517036, 517315, 517684, 518369, 518420, 518739, 520169, 520338, 520593, 521288, 521868, 522955, 524097, 525071, 525334, 525617, 527351, 527559, 528187, 529236, 529633, 530208, 530452, 531175, 531400, 532156, 533099, 533613, 533961, 534639, 535482, 535679, 535929, 536531, 536862, 537379, 537646, 537914, 538438, 539291, 539505, 539778, 541286, 542231, 542577, 542787, 543440, 544398, 544703, 545146, 545341, 545555, 547020, 547116, 547337, 547989, 548305, 548953, 549500, 552346, 553158, 554591, 555183, 557121, 557466, 557612, 558916, 559129, 559408, 559841, 560374, 560401, 560853, 561182, 561607, 561792, 562100, 563168, 563417, 564017, 564450, 564551, 566348, 566585, 567043, 567313, 567643, 568272, 568883, 570265, 570494, 570680, 572355, 572670, 572848, 574147, 574245, 575682, 575958, 576923, 578119, 578824, 579586, 579872, 580241, 580464, 580634, 581767, 582041, 582244, 583349, 583679, 583918, 584443, 584683, 584810, 585396, 585561, 587234, 587293, 587553, 588191, 588519, 588626, 588858, 589247, 589783, 592340, 592559, 592854, 594559, 594849, 595052, 596886, 597500, 597684, 598407, 598838, 599300, 599648, 600656, 600947, 602333, 603081, 603325, 603767, 603963, 604193, 605527, 606161, 606317, 606538, 607015, 607302, 607969, 608143, 608349, 608657, 608858, 609477, 610426, 610788, 611049, 611122, 611708, 612364, 613580, 614100, 614368, 614905, 615365, 617644, 618120, 619168, 619689, 619846, 620166, 621055, 621090, 622262, 622856, 624269, 624629, 625501, 625814, 626414, 627686, 627956, 629486, 629803, 630143, 630390, 631266, 631481, 632273, 632878, 633493, 633956, 634280, 635192, 635792, 636533, 637334, 637916, 638388, 638697, 638823, 639194, 639991, 640155, 641530, 642035, 642154, 642657, 643714, 644336, 644426, 644838, 645314, 646164, 646532, 646977, 647263, 647586, 648207, 648498, 649703, 650005, 650664, 650775, 651444, 651589, 652412, 652798, 652952, 653113, 653544, 654118, 654623, 654923, 655159, 655526, 656144, 656812, 657655, 658353, 658952, 659316, 659890, 661406, 661640, 662047, 662848, 663054, 663948, 664584, 664845, 665494, 666139, 666439, 666631, 667116, 667623, 668884, 669015, 670191, 670511, 671395, 671610, 671800, 672219, 672283, 672863, 674659, 675017, 676175, 676647, 677189, 677954, 678812, 680001, 680922, 680989, 681296, 681563, 683724, 683915, 684542, 684971, 685647, 686853, 688273, 688637, 688920, 690107, 693108, 694577, 695144, 695578, 695874, 696327, 696638, 696891, 697699, 698243, 698765, 699192, 699470, 700595, 700765, 701358, 702004, 703135, 703386, 703748, 704474, 705030, 705349, 706533, 706761, 707861, 710287, 710635, 711000, 712585, 713122, 714230, 714323, 716049, 716604, 716811, 717061, 717431, 717702, 717956, 718425, 718888, 719280, 719402, 719719, 720015, 720192, 720612, 720941, 721941, 722330, 724082, 724454, 724538, 724948, 725222, 725414, 726335, 728227, 728556, 728958, 729517, 729660, 730325, 731107, 731570, 731948, 732880, 732977, 733804, 734463, 734717, 734741, 735104, 735419, 735729, 736193, 736950, 737409, 737703, 737807, 738102, 738459, 738580, 739237, 739463, 739755, 740007, 740194, 740578, 741172, 741430, 741691, 742092, 742404, 743117, 743781, 744042, 745016, 745234, 746072, 746275, 746802, 747831, 748186, 748736, 749917, 750372, 750965, 751252, 752255, 752632, 753082, 753305, 753744, 754265, 754472, 755027, 755723, 757233, 757786, 758242, 758945, 759132, 759900, 761019, 761843, 762090, 762903, 763393, 764039, 764580, 764739, 765433, 767412, 767899, 768381, 768551, 769227, 769517, 769575, 769918, 770074, 770702, 771035, 771454, 771757, 771845, 772167, 772960, 773274, 774051, 774238, 774536, 776185, 776666, 776924, 777071, 778687, 778760, 779348, 779738, 779956, 780198, 780810, 781683, 781850, 782502, 782636, 783563, 784151, 784883, 786426, 786971, 788362, 788705, 789052, 789439, 789856, 790185, 791499, 792269, 792524, 792592, 794280, 794685, 795607, 795951, 796272, 796940, 798400, 799824, 800049, 802041, 802147, 802893, 803790, 803888, 804476, 805048, 806024, 806205, 806419, 807678, 807848, 808584, 808751, 809233, 809838, 810003, 810464, 810736, 811471, 811534, 811981, 812111, 812536, 813100, 814730, 816322, 816693, 816937, 817313, 818356, 818864, 819636, 819740, 820589, 821355, 821815, 822348, 822618, 822792, 823278, 824504, 824745, 825549, 826396, 826667, 827362, 827494, 827745, 828100, 828266, 828659, 829471, 829983, 830852, 831041, 831277, 831924, 833255, 834049, 835128, 835554, 835744, 836079, 836392, 837150, 838985, 839863, 840520, 841363, 842449, 842559, 843624, 844659, 845279, 847041, 847468, 847868, 847945, 848613, 849489, 850670, 850880, 851482, 851996, 852678, 852876, 853550, 854478, 855909, 856417, 857416, 857903, 858793, 859227, 859446, 860630, 861074, 861825, 862592, 862752, 863813, 864885, 865133, 865678, 865908, 866587, 866994, 867268, 867788, 867924, 868880, 869287, 869874, 869902, 871151, 871237, 871587, 871933, 872843, 873236, 873639, 873965, 874665, 875374, 876244, 876494, 876832, 877802, 878323, 878902, 879569, 880489, 881030, 881331, 881633, 882678, 883010, 883575, 884215, 884267, 885459, 885601, 886706, 887132, 887681, 888504, 888604, 889137, 890285, 890742, 891395, 891816, 893143, 893461, 895169, 896579, 896938, 897108, 898468, 898836, 899159, 899740, 899935, 900804, 901285, 901560, 901721, 902174, 903665, 903773, 905297, 905559, 906906, 909180, 909610, 910779, 911080, 911443, 911830, 911915, 912379, 912709, 913497, 913945, 914282, 914568, 915807, 916369, 916706, 917084, 917927, 918667, 918879, 919160, 919793, 919942, 920138, 920772, 921547, 922004, 922573, 923027, 924421, 925478, 926394, 926468, 927215, 927282, 927798, 928160, 928374, 929114, 929357, 929625, 929813, 930781, 930969, 931203, 931631, 934235, 934949, 935513, 936003, 936878, 937598, 938248, 938580, 939135, 939282, 940121, 940432, 940548, 941128, 941414, 941604, 941951, 942104, 942477, 942749, 943158, 944107, 944787, 946592, 947186, 947790, 948419, 948880, 949058, 949474, 949543, 949848, 950044, 950463, 951029, 951452, 951731, 952030, 952158, 952784, 952923, 953819, 954536, 955564, 955679, 955983, 956201, 957268, 958142, 958826, 959182, 959708, 960030, 960423, 960846, 962394, 962745, 963030, 963970, 964397, 964755, 966430, 966706, 967255, 967645, 967779, 968669, 969043, 969470, 970228, 971075, 971361, 972227, 972388, 973130, 973766, 974663, 975119, 975997, 976286, 978556, 978699, 978948, 979337, 979563, 981061, 981525, 982044, 982792, 983308, 983682, 984284, 984682, 985875, 986342, 986768, 987077, 987957, 988177, 988765, 989022, 989642, 991109, 991692, 992443, 992778, 993553, 994402, 994804, 995183, 996055, 996342, 996795, 996868, 997535, 997914, 998774, 999566, 1000019, 1000495, 1001670, 1001742, 1002131, 1002377, 1002678, 1003033, 1003684, 1004149, 1004375, 1004875, 1005149, 1005810, 1006164, 1007486, 1007672, 1007958, 1009048, 1009741, 1010029, 1010727, 1011659, 1012035, 1012337, 1012506, 1013568, 1013873, 1014398, 1014649, 1016702, 1017556, 1018275, 1018676, 1020086, 1020190, 1020544, 1020725, 1021142, 1021308, 1022007, 1022219, 1022648, 1022865, 1023866, 1024221, 1024459, 1024629, 1024960, 1025228, 1026565, 1028064, 1030393, 1030813, 1031001, 1031620, 1034217, 1034943, 1035336, 1035657, 1035920, 1036576, 1037072, 1037687, 1038558, 1039459, 1039732, 1040585, 1040873, 1040913, 1041854, 1042794, 1043382, 1043457, 1043824, 1044916, 1045442, 1045597, 1045805, 1046060, 1046519, 1046595, 1047574, 1047973, 1048203 );

  type key is array(0 to 63) of integer;
  constant answer_key : key :=
  ( 0, 1572882, 1310740, 3670035, 65564, 4128789, 1376268, 1310737, 7, 2490394, 1048598, 3932196, 1376276, 1114139, 2621464, 1376280, 8, 1048596, 2621474, 4128792, 7, 1, 1376267, 1310754, 2293771, 2883599, 14, 3670034, 31, 655383, 3670045, 1376270, 2031639, 1703959, 4128793, 1376265, 2621464, 1572887, 3014675, 983066, 2883600, 3866645, 2097182, 22, 4128777, 1310731, 524306, 458774, 3866644, 2818075, 3801109, 393258, 28, 393242, 13, 1572881, 2293773, 1703954, 65556, 4128784, 3538961, 1900572, 1638426, 8 );

  constant NUM_EDGES : integer := 1843;
  constant TEST_SIZE : integer := 64;
  constant MAX_CYCLES : integer  := TEST_SIZE*4;

  signal clk : std_logic := '0';
  signal rst : std_logic := '1';

  signal mmap_wr_en   : std_logic                         := '0';
  signal mmap_wr_addr : std_logic_vector(MMAP_ADDR_RANGE) := (others => '0');
  signal mmap_wr_data : std_logic_vector(MMAP_DATA_RANGE) := (others => '0');

  signal mmap_rd_en   : std_logic                         := '0';
  signal mmap_rd_addr : std_logic_vector(MMAP_ADDR_RANGE) := (others => '0');
  signal mmap_rd_data : std_logic_vector(MMAP_DATA_RANGE);

  signal sim_done : std_logic := '0';

begin

  UUT : entity work.user_app
    port map (
      clk          => clk,
      rst          => rst,
      mmap_wr_en   => mmap_wr_en,
      mmap_wr_addr => mmap_wr_addr,
      mmap_wr_data => mmap_wr_data,
      mmap_rd_en   => mmap_rd_en,
      mmap_rd_addr => mmap_rd_addr,
      mmap_rd_data => mmap_rd_data);

  -- toggle clock
  clk <= not clk after 5 ns when sim_done = '0' else clk;

  -- process to test different inputs
  process

    procedure clearMMAP is
    begin
      mmap_rd_en <= '0';
      mmap_wr_en <= '0';
    end clearMMAP;

    variable errors : integer := 0;

    variable result : std_logic_vector(C_MMAP_DATA_WIDTH-1 downto 0);
    variable done   : std_logic;
    variable count  : integer;

  begin
    report "============================SIMULATION START============================" severity note;
    -- reset circuit  
    rst <= '1';
    clearMMAP;
    wait for 200 ns;

    rst <= '0';
    wait until clk'event and clk = '1';
    wait until clk'event and clk = '1';

    -- write contents to input ram, which starts at addr 0
    --for i in 0 to (TEST_SIZE / 4) - 1 loop
    --  mmap_wr_addr <= C_MEM_IN_SEL_ADDR;
    --  mmap_wr_en   <= '1';
    --  mmap_wr_data <= std_logic_vector(to_unsigned(i, C_MMAP_DATA_WIDTH));
    --  wait until clk'event and clk = '1';
    --  clearMMAP;
    --  for j in 0 to TEST_SIZE - 1 loop
    --    mmap_wr_addr <= std_logic_vector(to_unsigned(j, C_MMAP_ADDR_WIDTH));
    --    mmap_wr_en   <= '1';
    --    mmap_wr_data <= std_logic_vector(to_unsigned(input_key(4*i, j), 8) &
    --                                     to_unsigned(input_key(4*i+1, j), 8) &
    --                                     to_unsigned(input_key(4*i+2, j), 8) &
    --                                     to_unsigned(input_key(4*i+3, j), 8));
    --    wait until clk'event and clk = '1';
    --    clearMMAP;
    --  end loop;      
    --end loop;

    --for i in 0 to TEST_SIZE - 1 loop
    --  mmap_wr_addr <= C_MEM_IN_SEL_ADDR;
    --  mmap_wr_en   <= '1';
    --  mmap_wr_data <= std_logic_vector(to_unsigned(i, C_MMAP_DATA_WIDTH));
    --  wait until clk'event and clk = '1';
    --  clearMMAP;
    --  for j in 0 to TEST_SIZE - 1 loop
    --    mmap_wr_addr <= std_logic_vector(to_unsigned(j, C_MMAP_ADDR_WIDTH));
    --    mmap_wr_en   <= '1';
    --    mmap_wr_data <= std_logic_vector(to_unsigned(input_key(i, j), 32));
    --    wait until clk'event and clk = '1';
    --    clearMMAP;
    --  end loop;      
    --end loop;

    for i in 0 to NUM_EDGES - 1 loop
     mmap_wr_addr <= std_logic_vector(to_unsigned(i, C_MMAP_ADDR_WIDTH));
     mmap_wr_en   <= '1';
     mmap_wr_data <= std_logic_vector(to_unsigned(edge_list(i), 32));
     wait until clk'event and clk = '1';
     clearMMAP;   
    end loop;   

    -- send size
    mmap_wr_addr <= C_SIZE_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(TEST_SIZE, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;

    -- send src
    mmap_wr_addr <= C_SRC_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(0, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;

    ---- send go = 1 over memory map
    mmap_wr_addr <= C_GO_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(1, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;
    
    done  := '0';
    count := 0;

    -- read the done signal every cycle to see if the circuit has
    -- completed.
    --
    -- equivalent to wait until (done = '1') for TIMEOUT;      
    while done = '0' and count < MAX_CYCLES loop

      mmap_rd_addr <= C_DONE_ADDR;
      mmap_rd_en   <= '1';
      wait until clk'event and clk = '1';
      clearMMAP;
      -- give entity one cycle to respond
      wait until clk'event and clk = '1';
      done         := mmap_rd_data(0);
      count        := count + 1;
    end loop;

    if (done /= '1') then
      errors := errors + 1;
      report "Done signal not asserted before timeout.";
    end if;

    -- read outputs from output memory
    for i in 0 to TEST_SIZE-1 loop
      mmap_rd_addr   <= std_logic_vector(to_unsigned(i, C_MMAP_ADDR_WIDTH));
      mmap_rd_en     <= '1';            
      wait until clk'event and clk = '1';
      clearMMAP;
      -- give entity one cycle to respond
      wait until clk'event and clk = '1';
      result := mmap_rd_data;

      if (unsigned(result) /= answer_key(i)) then
        errors := errors + 1;
        report "Result for " & integer'image(i) &
          " is incorrect. The output is " &
          integer'image(to_integer(unsigned(result))) &
          " but should be " & integer'image(answer_key(i));
      end if;
    end loop;  -- i

    report "SIMULATION FINISHED!!!";
    report "TOTAL ERRORS : " & integer'image(errors);
    report "=============================SIMULATION END=============================" severity note;
    sim_done <= '1';
    wait;

  end process;
end tb;
