../ip_repo/accelerator_1.0/src/mux_2_1.vhd