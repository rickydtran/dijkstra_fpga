-- Ricky Tran
-- University of Florida
-- user_app_tb.vhd

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.config_pkg.all;
use work.user_pkg.all;

entity user_app_tb is
end user_app_tb;

architecture tb of user_app_tb is
  type t_2d_a is array(0 to 63, 0 to 63) of integer range 0 to 255;
  constant input_key : t_2d_a :=
  ((    0,     0,     0,   211,     0,     0,     0,     0,     1,     0,     0,     0,     0,     0,     0,     0,     0,   175,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    58,     0,     0,     0,   106,     0,     0,     0,   127,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    70),
   (    0,     0,     0,     0,     0,     0,     0,    59,     0,     0,     0,     0,     0,     0,   191,     0,     0,     0,     0,     0,   130,     0,   154,     0,     0,     0,     0,     0,   183,     0,     0,     0,     0,     0,     0,     0,     0,     0,     9,     0,     0,     0,     0,     0,   217,     0,     0,     0,    71,     0,     0,     0,     0,     0,     0,     0,     0,   147,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,   141,     0,     0,     0,     0,   239,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   239,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (  211,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   250,    55,    15,     0,     0,     0,     0,     0,    73,     0,     0,     0,     0,     0,   242,     0,     0,    70,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,   141,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   160,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   239,   231,     0,     0,   166,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   175,     0,     0,     0,     0,     0,     0,   244,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   138,     0,     0,     0,     0,     0,     0,     0,   236,     0,   245,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    26),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,   160,     0,   190,     0,     0,     0,     0,     0,     0,     0,    51,     0,     0,    17,     0,    34,     0,     0,     0,     0,     0,     0,     0,   213,   134,   192,     0,   231,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   101,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,    59,     0,     0,     0,     0,     0,     0,     0,     0,    72,     0,     0,     0,     0,     0,   186,     0,     0,     6,     0,     0,     0,     0,     0,   165,   146,     0,     0,     0,     0,     0,     3,     0,     0,     0,     0,     0,     0,     0,   136,   127,     0,     0,     0,    16,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    94,     0,     0),
   (    1,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   183,     0,    13,     0,     0,     0,     0,     0,     0,     0,     0,     0,    96,     0,     0,   130,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   119,     0,     0,   173,     0,     0,     0,     0),
   (    0,     0,   239,     0,     0,     0,   160,     0,     0,     0,     0,     0,     0,     0,     0,   172,     0,     0,     0,     0,   158,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   210,     0,     0,     0,   107,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    42),
   (    0,     0,     0,     0,     0,     0,     0,    72,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    45,    36,     0,     0,   124,     0,     0,     0,     0,     0,     0,    94,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    28,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,   190,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   193,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,   183,     0,     0,     0,     0,     0,     0,   131,     0,     0,     0,     0,    61,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   255,     0,     0,     0,     0,     0,     0,     0,   226,     0,     0,     0,     0,     0,     0,     0,     0,     0,    29,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   249,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   165,     0,     0,     0,     0,     0,     0,     0,     0,     0,   140,     0,     0,     0,     0,     0,     0,     0,   227,     0,     0,     0,     0,     0,     0,   170,     0,     0,     0),
   (    0,   191,     0,     0,     0,     0,     0,     0,    13,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   215,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   207,     0,   213,    86,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   120,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,   172,     0,     0,   131,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    58,   147,   134,     0,     0,     0,     0,     9,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   229,   132,     0,     0,     0,     0,     0,     0,    31,     0,     0,     0,     0,    67,     0,    62,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,   186,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   158,     0,     0,     0,     0,     0,     0,     0,     0,     0,    44,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (  175,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    40,     0,     0,     0,     0,     0,     0,     0,   205,    89,     0,     0,     0,     0,     0,     0,     0,     0,   244,     0,     0,     0,   131,     0,     0,     0,   229,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    19,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   224,    87,     0,     0,     0,    69,     0,     0,     0,   247,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,    51,     6,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   197,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,   130,     0,     0,     0,   175,     0,     0,     0,   158,     0,     0,    61,     0,   215,     0,   158,     0,     0,     0,     0,     0,     0,    87,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   196,     0,     0,     0,     0,     0,     0,   227,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    92,     0,     0,     0,     0,     0,   118,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    71,     0,   126,     0,     0,     0,     0,     0),
   (    0,   154,     0,   250,   160,     0,    17,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    40,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   243,     0,   240,   216,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   106),
   (    0,     0,     0,    55,     0,     0,     0,     0,     0,     0,    45,     0,     0,   249,     0,    58,     0,     0,     0,     0,    87,    92,     0,     0,     0,   117,     0,     0,     0,     0,    55,     0,     0,     0,     0,     0,     0,     0,     0,   228,     0,    25,     0,     0,   157,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   159,     0,     0),
   (    0,     0,     0,    15,     0,     0,    34,     0,    96,     0,    36,     0,     0,     0,     0,   147,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    97,     0,    13,     0,    86,     0,     0,     0,     0,     0,     0,     0,   252,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   172,     0,     0,     0,    89,     0,     0,     0,   217),
   (    0,     0,     0,     0,     0,     0,     0,   165,     0,     0,     0,     0,     0,     0,     0,   134,     0,     0,     0,     0,     0,     0,     0,   117,     0,     0,     0,     0,     0,     0,     0,     0,     0,   179,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     3,    33,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,   146,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   175,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     6,   152,   116,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,   244,     0,     0,   130,     0,   124,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   186,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    72,     0,    46,     0,     0,     0,   143,    48,   248,     0,     0,    55,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,   183,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    19,     0,     0,     0,     0,     0,     0,     0,     0,   186,     0,     0,   161,     0,     0,     0,   238,     0,     0,   253,   188,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   177,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   118,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   129,     0,     0,     0,     0,     0,     0,     0,   160,     0,     0,     0,     0,   218,     0,   220,     0,     0,     0,     0,     0),
   (    0,     0,     0,    73,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     9,    44,   205,     0,     0,     0,     0,     0,    55,     0,     0,     0,     0,   161,     0,     0,    28,   112,     0,     0,     0,     0,   178,     0,     0,     0,     0,     0,     0,     0,     0,   193,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    89,     0,     0,     0,     0,     0,     0,    97,     0,     0,     0,     0,     0,    28,     0,     0,     0,     0,     0,     0,     0,     0,    56,     0,     0,     0,   102,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,   213,     3,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   112,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    35,     0,   150,     0,     0,   148,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (   58,     0,     0,     0,     0,     0,   134,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    13,   179,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   249,     0,     0,     0,     0,     0,     0,     0,   125,     0,     0,   158,     0,   247,     0,     0,   245,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,   192,     0,     0,     0,    94,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   238,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    41,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   165,   207,     0,     0,     0,     0,     0,     0,     0,     0,     0,    86,     0,   175,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   241,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   154,     0,     0,    57,     0),
   (    0,     0,     0,   242,     0,     0,   231,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (  106,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   213,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   253,     0,   178,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   245,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     9,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    86,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   188,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    66,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,    70,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   196,     0,     0,   228,     0,     0,     0,     0,     0,     0,     0,    56,     0,     0,     0,     0,     0,     0,     0,     0,     0,   231,     0,   127,     0,     0,   255,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,   136,     0,     0,     0,     0,     0,     0,     0,     0,     0,   244,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    23,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (  127,     0,     0,     0,     0,     0,     0,   127,     0,     0,     0,     0,   255,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    25,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   241,     0,     0,     0,   231,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   190,     0,     0,     0,     0,     0,     0,     0,   144,     0,     0,     0),
   (    0,     0,     0,     0,     0,   138,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   224,   197,     0,     0,     0,     0,     0,     0,     0,    72,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    23,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   214,     0,     0,     0,     0,     0,     0,     0,     0,     0,    11,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    87,     0,     0,     0,     0,     0,   252,     0,     0,     0,     0,   129,     0,   102,     0,     0,     0,     0,     0,     0,     0,   127,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    38,     0,   116,     0,     0,     0,     0,     0,     0,     0,     0,    58,    35,     0),
   (    0,   217,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   131,     0,     0,     0,     0,     0,   157,     0,     0,     0,    46,     0,     0,     0,     0,     0,   249,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   127,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,   239,     0,     0,    16,     0,     0,     0,     0,     0,   140,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    35,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,   239,     0,   231,     0,     0,     0,     0,   210,     0,     0,     0,     0,     0,   229,     0,     0,     0,     0,   227,     0,     0,     0,     0,     0,     0,     0,     0,     0,   193,     0,     0,     0,     0,     0,     0,     0,     0,   255,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   132,     0,     0,    69,     0,     0,     0,   243,     0,     0,     0,     0,     0,     0,     0,     0,     0,   150,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   129,     0,     0,   251,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,    71,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   229,     0,     0,     0,     0,     0,     0,     0,     0,     0,   143,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    66,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   182,     0,     0),
   (    0,     0,     0,     0,   166,     0,     0,     0,     0,     0,     0,     0,   226,     0,   120,     0,     0,     0,     0,     0,     0,     0,   240,     0,     0,     0,     0,    48,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   129,     0,     0,     0,     0,   139,     0,     0,     0,     0,     0,     0,     0,   185,     0,     0,     0),
   (    0,     0,     0,     0,     0,   236,     0,     0,     0,   107,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   216,     0,     0,     0,     0,   248,     0,     0,     0,     0,   148,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    38,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   247,     0,     0,     0,     0,     0,     0,     0,     6,     0,     0,   160,     0,     0,     0,     0,    41,     0,     0,   245,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   193,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,   245,     0,     0,     0,     0,    28,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   152,     0,     0,     0,     0,     0,     0,   125,     0,     0,     0,     0,     0,     0,     0,   190,   214,   116,     0,     0,     0,   251,     0,   139,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   248,     0),
   (    0,     0,     0,     0,     0,     0,   101,     0,     0,     0,     0,     0,     0,   227,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     3,   116,    55,   177,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   127,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   210,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    31,     0,     0,     0,     0,     0,     0,     0,     0,     0,    33,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    77,   198,     0,     0,    51,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   172,     0,     0,     0,     0,     0,     0,     0,     0,   158,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    77,     0,   169,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,   119,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    71,     0,     0,     0,     0,     0,     0,     0,   218,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   198,   169,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,   147,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   247,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   210,     0,     0,     0,     0,   244,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   126,     0,     0,     0,     0,     0,     0,     0,   220,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   193,     0,     0,     0,     0,     0,   244,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,   173,     0,     0,   193,    29,     0,     0,    67,     0,     0,     0,     0,     0,     0,     0,     0,    89,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   154,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    51,     0,     0,     0,     0,     0,     0,     0,    64,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   170,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   245,     0,     0,     0,     0,     0,     0,     0,   144,     0,     0,     0,     0,     0,     0,     0,   185,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,    94,     0,     0,     0,     0,     0,     0,     0,    62,     0,     0,     0,     0,     0,     0,     0,   159,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    58,     0,     0,     0,     0,   182,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0),
   (    0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,    57,     0,     0,     0,     0,     0,     0,    11,    35,     0,     0,     0,     0,     0,     0,     0,     0,   248,     0,     0,     0,     0,     0,     0,    64,     0,     0,     0,   205),
   (   70,     0,     0,     0,     0,    26,     0,     0,     0,    42,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   106,     0,   217,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,     0,   205,     0));
   
  type key is array(0 to 63) of integer;
  constant answer_key : key :=
  ( 0, 2490477, 590175, 1572950, 1442074, 4128864, 1572969, 1245346, 1, 4128880, 1572971, 393511, 524472, 2949438, 524302, 1966248, 1966283, 1441954, 1835315, 393372, 1507556, 3670207, 393338, 196749, 2162759, 3473597, 3342584, 524419, 2490656, 1376565, 196767, 1573032, 458917, 58, 655561, 1573021, 196936, 106, 917604, 196764, 2752738, 127, 1769675, 4063481, 1769649, 458930, 590146, 3211527, 2490534, 917638, 590043, 2228466, 655495, 1769658, 983239, 2162904, 524408, 65792, 1376573, 1573024, 2687247, 983270, 2293974, 70 );

  constant TEST_SIZE : integer := 64;
  constant MAX_CYCLES : integer  := TEST_SIZE*4;

  signal clk : std_logic := '0';
  signal rst : std_logic := '1';

  signal mmap_wr_en   : std_logic                         := '0';
  signal mmap_wr_addr : std_logic_vector(MMAP_ADDR_RANGE) := (others => '0');
  signal mmap_wr_data : std_logic_vector(MMAP_DATA_RANGE) := (others => '0');

  signal mmap_rd_en   : std_logic                         := '0';
  signal mmap_rd_addr : std_logic_vector(MMAP_ADDR_RANGE) := (others => '0');
  signal mmap_rd_data : std_logic_vector(MMAP_DATA_RANGE);

  signal sim_done : std_logic := '0';

begin

  UUT : entity work.user_app
    port map (
      clk          => clk,
      rst          => rst,
      mmap_wr_en   => mmap_wr_en,
      mmap_wr_addr => mmap_wr_addr,
      mmap_wr_data => mmap_wr_data,
      mmap_rd_en   => mmap_rd_en,
      mmap_rd_addr => mmap_rd_addr,
      mmap_rd_data => mmap_rd_data);

  -- toggle clock
  clk <= not clk after 5 ns when sim_done = '0' else clk;

  -- process to test different inputs
  process

    procedure clearMMAP is
    begin
      mmap_rd_en <= '0';
      mmap_wr_en <= '0';
    end clearMMAP;

    variable errors : integer := 0;

    variable result : std_logic_vector(C_MMAP_DATA_WIDTH-1 downto 0);
    variable done   : std_logic;
    variable count  : integer;

  begin
    report "============================SIMULATION START============================" severity note;
    -- reset circuit  
    rst <= '1';
    clearMMAP;
    wait for 200 ns;

    rst <= '0';
    wait until clk'event and clk = '1';
    wait until clk'event and clk = '1';

    -- write contents to input ram, which starts at addr 0
    for i in 0 to (TEST_SIZE / 4) - 1 loop
      mmap_wr_addr <= C_MEM_IN_SEL_ADDR;
      mmap_wr_en   <= '1';
      mmap_wr_data <= std_logic_vector(to_unsigned(i, C_MMAP_DATA_WIDTH));
      wait until clk'event and clk = '1';
      clearMMAP;
      for j in 0 to TEST_SIZE - 1 loop
        mmap_wr_addr <= std_logic_vector(to_unsigned(j, C_MMAP_ADDR_WIDTH));
        mmap_wr_en   <= '1';
        mmap_wr_data <= std_logic_vector(to_unsigned(input_key(4*i, j), 8) &
                                         to_unsigned(input_key(4*i+1, j), 8) &
                                         to_unsigned(input_key(4*i+2, j), 8) &
                                         to_unsigned(input_key(4*i+3, j), 8));
        wait until clk'event and clk = '1';
        clearMMAP;
      end loop;      
    end loop;

    -- send size
    mmap_wr_addr <= C_SIZE_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(TEST_SIZE, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;

    -- send src
    mmap_wr_addr <= C_SRC_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(0, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;

    ---- send go = 1 over memory map
    mmap_wr_addr <= C_GO_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(1, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;
    
    done  := '0';
    count := 0;

    -- read the done signal every cycle to see if the circuit has
    -- completed.
    --
    -- equivalent to wait until (done = '1') for TIMEOUT;      
    while done = '0' and count < MAX_CYCLES loop

      mmap_rd_addr <= C_DONE_ADDR;
      mmap_rd_en   <= '1';
      wait until clk'event and clk = '1';
      clearMMAP;
      -- give entity one cycle to respond
      wait until clk'event and clk = '1';
      done         := mmap_rd_data(0);
      count        := count + 1;
    end loop;

    if (done /= '1') then
      errors := errors + 1;
      report "Done signal not asserted before timeout.";
    end if;

    -- read outputs from output memory
    for i in 0 to TEST_SIZE-1 loop
      mmap_rd_addr   <= std_logic_vector(to_unsigned(i, C_MMAP_ADDR_WIDTH));
      mmap_rd_en     <= '1';            
      wait until clk'event and clk = '1';
      clearMMAP;
      -- give entity one cycle to respond
      wait until clk'event and clk = '1';
      result := mmap_rd_data;

      if (unsigned(result) /= answer_key(i)) then
        errors := errors + 1;
        report "Result for " & integer'image(i) &
          " is incorrect. The output is " &
          integer'image(to_integer(unsigned(result))) &
          " but should be " & integer'image(answer_key(i));
      end if;
    end loop;  -- i

    report "SIMULATION FINISHED!!!";
    report "TOTAL ERRORS : " & integer'image(errors);
    report "=============================SIMULATION END=============================" severity note;
    sim_done <= '1';
    wait;

  end process;
end tb;
