../ip_repo/accelerator_1.0/src/decoder_edge.vhd