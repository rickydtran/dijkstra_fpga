../ip_repo/accelerator_1.0/src/comp_min.vhd