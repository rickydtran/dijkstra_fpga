-- Ricky Tran
-- University of Florida
-- user_app_tb.vhd

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.config_pkg.all;
use work.user_pkg.all;

entity user_app_tb is
end user_app_tb;

architecture tb of user_app_tb is
  type t_2d_a is array(0 to 127, 0 to 127) of integer range 0 to 255;
  constant input_key : t_2d_a :=
  ((    0,    95,    88,   174,     5,   177,   192,     5,     0,     0,    70,    57,   238,   190,     0,   109,   135,   166,   123,   174,    42,     8,   171,     1,   213,     0,   142,   131,     0,   184,    80,    98,   124,   139,   146,    47,   220,     0,   129,   198,    63,    36,   117,   219,    38,   198,   212,   184,    29,   123,   248,   192,   224,   172,     7,   130,     7,    68,    97,   198,    77,    49,   175,   202,     8,    39,   240,   185,   126,   131,    33,    62,   150,    96,   248,   102,   105,   245,    74,    25,   138,    55,    27,   160,    11,   128,   162,   111,    15,    39,   242,    41,   212,   139,   225,    48,   173,   205,   179,   153,    89,    87,    49,     0,   181,   208,   137,   157,    92,   234,     0,   113,     0,   113,    56,   170,   248,   249,    47,   210,   114,    46,   127,   207,    57,    33,   139,   214),
   (   95,     0,   207,    13,     0,   114,   174,     0,   211,   179,    28,    86,   198,    51,     2,     0,   188,    27,   106,   137,   146,    17,    45,   126,   213,    60,   217,     0,   203,    55,   125,   202,   209,   251,    48,   171,    95,    57,   101,   214,   155,    57,    82,   173,   169,     0,   170,    64,    42,   135,     0,    29,   234,    83,   165,   127,   237,    43,     0,    35,   113,   253,    48,    53,    53,     0,   239,     3,    64,    90,    40,    30,   244,    37,    24,   105,     0,   213,   200,   182,   103,   234,     0,   232,   214,    43,   193,   118,    51,   235,    70,   110,    62,    51,    13,    36,    90,    46,   190,    38,   104,   152,   100,   248,   143,   236,   243,   137,    71,   191,    90,   191,   228,   174,    83,   163,    45,     1,     2,   166,    35,   250,    99,   137,    86,    32,   214,   240),
   (   88,   207,     0,   192,   167,   113,   142,     3,   237,   128,    26,    93,   104,   121,    15,     7,    44,   103,    42,   186,   118,   145,    99,   253,    23,   208,   178,    18,    99,   166,   202,   248,     2,   170,    59,   140,   220,   212,    93,     3,    77,   142,    46,   186,     0,   230,    24,    48,   232,   205,    70,   239,   118,    29,   140,   175,   165,    43,   249,   196,   250,     4,    52,    73,   179,    63,   187,    18,    37,    36,     0,    82,    46,   136,   197,   124,   196,    89,   181,     0,    75,   178,    14,   216,   244,    83,   150,   131,   114,   206,     0,   150,   218,     0,   200,     0,   251,   111,   195,   247,     0,    49,   209,   140,   189,   156,    88,    51,   132,     0,   232,    23,    68,   194,   252,    56,   193,   122,     0,    54,   169,    62,   218,   172,    70,    11,   137,    97),
   (  174,    13,   192,     0,     0,    82,    76,    73,   185,   233,   138,    41,   195,   168,   139,   170,    25,   137,   181,    49,    53,   209,    75,   116,     1,   103,   110,    87,   141,   201,   239,    81,   246,     0,   230,   119,   166,     0,    75,   204,    25,   213,    78,    75,   122,    68,    38,     0,    33,   249,   231,    76,   157,    41,   204,   214,   213,   121,   141,    42,    75,    67,     0,   229,   183,    16,   157,   184,   113,   122,    80,   131,   177,     0,    62,   190,     3,    38,    63,   147,     0,   125,   199,   182,   107,   241,   159,    77,   179,     0,   155,   135,    18,     0,   197,   135,    88,   149,    40,   188,    31,   153,    72,   131,   131,     0,   247,    43,   114,   218,    88,    15,   138,   160,   145,   125,   143,    41,   246,    76,   113,   152,    43,   160,    72,   169,    48,   105),
   (    5,     0,   167,     0,     0,   109,   199,   225,    67,   201,   153,   175,   156,   246,   183,   196,     0,    47,   165,    34,    25,    80,     5,    77,   253,   197,    94,   220,    57,   156,    61,    39,    60,    37,   248,   183,    15,    86,   117,    68,   207,    77,    25,    71,   109,     0,   146,   149,    25,   210,   253,   102,     4,   110,   233,     1,    68,   181,   117,   168,    88,   164,   248,   129,   192,   175,   142,   122,    70,     0,   147,   161,   111,   146,   203,    51,   142,    46,     0,     0,    19,   240,   238,   104,     0,   194,    23,   232,   215,     6,   180,   197,     0,   134,   207,   179,     0,   186,   132,   166,   233,     0,   223,   244,     0,    83,   199,   228,   125,   194,   222,   158,    80,    68,    76,     0,   237,    61,   196,   215,   111,   148,    44,    73,     0,   101,     0,   254),
   (  177,   114,   113,    82,   109,     0,    17,   110,   248,    33,    13,   130,    70,     3,   194,    95,   210,   101,   232,    71,     0,   184,    91,   133,   229,    88,    52,   161,   191,     0,   162,   159,   242,     0,    66,    64,    63,   213,   218,   147,   198,   105,    44,    17,   204,    64,   114,   211,    69,    49,   137,   156,   236,   181,     0,   161,    30,     0,   172,   127,   184,    66,   125,    91,     0,    33,    72,    21,   250,   175,    79,   197,     0,   228,   250,   217,    51,   167,    95,    18,   226,    28,   117,    15,     0,   196,   112,   246,   127,   105,   139,   214,    97,   216,     0,   190,    93,     0,     0,    36,   178,   143,    25,   116,   226,   136,   206,   229,   227,   229,    69,    86,    29,   111,   133,   167,    86,   122,    74,   122,   206,    53,   190,   146,     0,     7,   255,     0),
   (  192,   174,   142,    76,   199,    17,     0,     0,   244,   172,     0,    50,    95,    21,   211,   174,    96,    98,   187,    42,   169,    23,    62,   212,   114,   100,    16,    28,   190,    39,   145,   218,    69,    60,   183,     0,    60,   211,     0,    98,   197,   108,   132,     9,   147,     0,   166,     5,    81,   230,    18,   184,    55,   199,   131,   167,   183,   143,   173,     0,   173,    33,   117,    15,    13,   248,   201,   168,    29,     0,     0,   131,    97,   193,    83,     5,   184,   247,    35,   183,   233,   134,   132,     0,    80,     2,   228,   161,     0,   235,    16,   214,     6,   148,   219,    31,   168,    45,   223,   190,   201,    92,   134,   245,    33,   238,   225,   188,   186,   189,     0,     0,   164,    32,    34,   125,     0,   183,   191,    45,   182,    40,    79,   141,     3,   253,   212,   192),
   (    5,     0,     3,    73,   225,   110,     0,     0,   177,   201,   131,   142,   181,   154,     0,     0,   177,   132,   234,    57,    78,   132,    11,     0,    71,    79,   108,     1,   204,   136,   145,     5,   232,    19,    31,    55,    42,   137,     0,    80,    75,   202,     0,   206,   193,   253,   169,    11,    30,   231,    70,     4,     0,    51,     2,   129,   235,    70,    39,    88,     0,   243,    97,     7,   153,   191,   101,    47,   219,     0,    57,   156,   106,   205,    54,    56,    76,   140,   215,   182,   155,   105,   251,   105,    30,   112,   252,     0,     0,   159,     0,   182,   208,     2,    52,   192,   193,    43,    46,   107,    62,    99,    50,   174,    19,   216,   164,   117,   118,   219,     0,    10,   214,    26,    21,    81,    66,    91,    95,    67,   202,     0,   127,   141,   249,   182,   132,    61),
   (    0,   211,   237,   185,    67,   248,   244,   177,     0,   198,    42,    71,   199,   139,   205,   100,    84,    68,   171,   146,   151,     0,    95,   147,    62,   100,   109,   251,   255,    47,    21,   232,   250,     0,    22,   137,   171,    51,   122,    66,   142,    52,    82,   186,   132,   201,   223,    91,     0,   201,   150,     0,   236,   252,   179,   216,   163,    57,   191,   134,     0,   223,   197,   186,   123,   133,   113,   157,    58,    65,    66,   232,   105,   104,   177,    70,     0,    47,   183,    10,   139,     0,    57,   137,   155,   150,   189,   224,   208,   112,    86,   107,   199,    26,    48,   151,     9,    90,   209,   113,     0,    81,   135,   108,    86,     0,   233,    54,     0,    29,    52,   242,   159,   139,    17,   217,    24,   110,    36,   167,   126,   138,    72,   232,   102,   223,    59,    80),
   (    0,   179,   128,   233,   201,    33,   172,   201,   198,     0,    89,   150,    79,     0,    90,    52,   158,   162,    57,     0,   148,     0,   248,     0,    66,    73,   166,   225,    79,   152,   233,     0,    92,    66,     0,    48,     0,   142,    24,     0,   219,   135,   240,   214,   219,   107,   103,   217,   252,   236,   159,    94,   146,    44,   169,    25,    48,    96,   109,   158,    95,    14,   196,    92,    77,    43,   178,   247,   123,   159,   172,   104,   160,     0,   162,   101,   188,    95,    23,     0,   113,   241,   231,   128,    27,   253,   189,   176,    11,   127,    13,    63,    53,    41,    72,   115,   104,   153,    95,   169,   246,   134,    52,   159,    88,     0,    31,   188,     0,   214,    16,   123,   117,    33,    88,   244,   121,   167,    27,    24,    46,    16,   132,    19,   120,   153,    25,   249),
   (   70,    28,    26,   138,   153,    13,     0,   131,    42,    89,     0,    13,    78,   205,   238,   125,    60,    36,   200,   143,    64,    33,    85,   121,    15,   139,    36,   144,   133,     0,   135,     0,   208,    28,   117,    70,   110,   247,    81,    94,   191,   252,   233,   148,   159,     0,   107,    34,    15,    67,   157,   149,     0,    43,   245,     0,   131,   195,     0,    43,   143,    62,    27,   157,   142,   255,    46,   248,   251,    61,   197,    25,   141,    18,   253,   142,    19,   121,    68,   176,    15,     3,    76,     0,    91,   114,    96,     5,   154,    64,    51,    61,   150,    32,    93,   162,   172,   230,   110,   136,    58,    98,     0,   242,    70,    94,     7,     0,    93,   197,     0,   122,    24,   168,   156,    94,   248,   137,   190,   116,   146,    97,   120,     0,    48,    34,    54,     0),
   (   57,    86,    93,    41,   175,   130,    50,   142,    71,   150,    13,     0,    67,   234,   107,   133,   103,   209,    81,     0,   194,   129,    34,   195,    48,   215,    93,     3,   135,   201,   167,    71,     1,   156,   184,   153,   189,    70,    54,   199,     0,   202,   105,    25,   206,    89,    57,     0,   130,   152,    25,     0,   181,   111,   252,     0,    74,   222,   159,   199,    92,   244,    50,   244,   145,    20,   153,     7,    26,   133,   177,    51,   152,   125,   135,     0,   201,   206,    68,   132,    64,   204,   162,   143,   178,   111,   185,   227,   146,    65,    75,   187,   152,   194,    73,   126,   173,    72,   252,   180,   185,   201,   132,    39,   207,   221,   175,   255,     0,    52,   133,   107,    96,   130,   111,   178,   187,    99,   122,    50,    43,   216,    20,   229,     1,   146,   173,   195),
   (  238,   198,   104,   195,   156,    70,    95,   181,   199,    79,    78,    67,     0,    90,    75,    43,    35,   148,     0,   179,    50,   245,   133,   156,    66,   109,    49,   154,    66,   100,   231,    47,   141,    21,    40,     9,    13,   225,   116,    93,   145,   155,   247,   214,     8,   158,     0,    90,    50,   162,    59,   190,   129,    73,   137,    88,    60,   107,   170,     0,     0,   163,    59,   104,    46,    97,   135,    95,     0,    87,   177,    85,    15,    52,   204,   155,   237,    63,   102,    72,   176,   140,   227,    53,     0,   151,    46,   177,    27,   181,   115,    25,   138,   123,    57,    16,   190,    36,   213,    58,    99,   106,    65,   153,   209,   196,   146,   253,   147,   168,    69,     2,   136,   161,   254,   141,   161,    27,   224,     0,   219,     0,   213,   103,    97,    60,     0,     0),
   (  190,    51,   121,   168,   246,     3,    21,   154,   139,     0,   205,   234,    90,     0,    87,     0,   142,   204,    58,   172,   121,   183,    67,   252,    82,   158,   239,   177,   119,    74,   188,   158,   139,     0,    76,    91,   211,   173,   240,    13,    70,   182,   195,     0,    98,   121,     5,   117,   134,   159,   143,    73,    69,    61,    25,   162,   130,    63,    23,   133,   118,   175,   115,   208,   204,    84,     0,   223,   251,    34,   186,   171,     0,   164,   110,   100,     0,   253,   192,     2,    94,   176,     0,   114,    56,   225,     0,    88,    72,     0,   208,    78,   248,    99,   175,    33,   204,   190,   130,    97,   100,   244,    43,   107,    93,   171,   109,   156,   193,   137,    24,     0,   197,     2,   252,    25,    47,   187,   128,    54,   147,   103,   100,   165,   156,   214,    72,    33),
   (    0,     2,    15,   139,   183,   194,   211,     0,   205,    90,   238,   107,    75,    87,     0,   213,   238,    65,   132,   229,   131,   177,   152,    78,   183,   118,    26,    87,   158,    96,    24,    39,   204,    83,     0,   123,   156,    24,    90,   234,   209,     0,    93,   104,    22,    47,   246,   189,   236,   149,   237,   224,     0,    32,   111,   254,   228,   152,   196,    60,   125,    96,    98,    93,    36,   239,    76,   159,   110,   203,   140,    37,    58,   108,     0,    62,   198,    52,   250,    25,    31,    71,     0,   228,   134,    33,   190,   167,    19,   188,   177,    41,     1,   153,     0,     4,   235,   151,   200,     0,    79,   145,    29,   186,   231,   164,   247,   151,    19,   159,    19,    46,    37,    97,    19,    91,   214,   199,   130,    14,    20,   156,    11,   186,    38,     0,    95,   125),
   (  109,     0,     7,   170,   196,    95,   174,     0,   100,    52,   125,   133,    43,     0,   213,     0,    17,   135,    56,   214,    42,    37,    13,    60,   144,   140,    83,   157,   219,   210,   112,   168,    62,    47,   211,   185,   244,   231,   130,    66,   151,   168,     0,   149,   200,   210,   184,   178,    94,   141,    83,   100,   209,   155,   100,    48,   110,    16,   184,   164,   187,   201,   129,   146,   233,    17,    50,    23,   235,    42,    94,   150,   141,   174,    79,     0,   214,   114,   234,   136,    93,    30,    59,   206,    46,   232,   147,    24,   171,    56,   236,    32,     9,   199,   144,   218,   163,   236,   209,    60,   101,   153,    75,    86,   151,   202,   172,   126,     8,    57,   192,    66,    54,    34,   227,     0,   243,    65,    85,   232,   235,   108,     0,   206,   194,     0,    56,   130),
   (  135,   188,    44,    25,     0,   210,    96,   177,    84,   158,    60,   103,    35,   142,   238,    17,     0,   252,   193,    34,   180,   114,   220,    44,   115,   118,   191,    64,   115,    63,   201,   100,   145,   102,   103,   194,   166,     0,   202,   226,   198,     0,   101,    82,    51,   183,    79,    18,   162,   137,    98,   157,    80,    63,    92,   168,     0,    52,   174,   102,   167,   160,    94,   221,   179,    41,    22,   230,    49,   112,   122,   113,    40,   119,     0,   158,   168,    25,   126,    91,     0,   212,   174,    47,    65,   254,   146,   138,   133,    12,   211,   113,   216,   220,   137,   254,    18,   210,   208,   237,    46,   188,   136,     0,   233,    38,    72,    39,    83,   202,    62,    51,   182,     0,    15,   234,   179,   217,   252,   145,   131,   175,    44,     1,   137,   169,     0,   134),
   (  166,    27,   103,   137,    47,   101,    98,   132,    68,   162,    36,   209,   148,   204,    65,   135,   252,     0,   177,   157,   166,   115,   236,   134,   103,    91,   215,   182,     0,   191,    82,    11,   213,   192,    25,   141,   221,   200,   155,   237,   222,   152,     0,   223,   120,   193,   210,    44,     0,    94,   112,    96,   197,   157,    27,   177,    52,   222,    34,   164,   180,    60,   124,    68,    11,    41,    78,   138,     2,    99,    86,   106,   102,   122,   179,     0,   233,    92,     0,    22,     5,   127,   153,     0,   105,   254,     0,   202,   111,   179,   132,   224,   105,   119,     4,   124,   210,   175,    52,    11,   143,   202,    87,    99,    47,   184,   141,   170,    22,    87,   214,   225,    62,    69,    83,   211,    27,   167,    75,    86,   108,    70,   151,     0,   131,   110,    52,   162),
   (  123,   106,    42,   181,   165,   232,   187,   234,   171,    57,   200,    81,     0,    58,   132,    56,   193,   177,     0,   168,    96,     7,   193,   103,   108,   196,    54,    39,   135,     0,   123,   162,    77,   180,    56,    19,   148,    14,    82,    78,    59,   101,    10,     0,   186,   210,    96,     0,     0,     0,   167,   168,   187,     1,    65,   206,     0,     5,    33,     0,    90,    10,   187,   250,   173,   254,    77,   122,     1,   165,   192,   238,   213,   175,   111,   241,     0,    39,   243,     0,   252,    48,   165,    62,    53,     0,   179,     0,   105,    24,   229,   174,    24,    94,    13,   189,    10,     0,    46,    14,   213,   249,    39,     0,    24,   197,     8,   189,   103,   234,   255,   159,     8,   185,     0,    35,   136,    40,    32,    70,    18,   211,   242,   165,    24,     0,   152,    72),
   (  174,   137,   186,    49,    34,    71,    42,    57,   146,     0,   143,     0,   179,   172,   229,   214,    34,   157,   168,     0,    23,    18,   168,    97,     0,    97,    98,     0,    95,    70,    66,   181,   104,     6,    95,   242,   106,   129,     0,    19,    26,    71,    22,   182,    72,    15,    37,    83,    24,    84,   137,     1,    21,   131,   179,    67,   166,   149,    58,   180,   235,    78,     0,    48,    27,    85,   126,    30,   173,   150,     2,    50,   110,   183,   110,   249,   173,    95,   227,    63,    32,   195,   211,   124,    65,    62,    63,   218,   180,    13,   248,    93,   209,   178,     0,     0,    14,   110,   141,    96,    73,    54,   150,   173,   242,    95,    44,    64,   112,     0,   248,    27,     0,    46,   254,   103,     5,    47,   102,   109,   137,   157,    45,   195,    67,     6,    64,   253),
   (   42,   146,   118,    53,    25,     0,   169,    78,   151,   148,    64,   194,    50,   121,   131,    42,   180,   166,    96,    23,     0,   190,   146,   181,   130,   213,   176,   253,   216,   218,   234,   153,   252,   120,   202,   161,   245,    78,    81,    65,   225,   212,    86,     0,   152,   231,   123,    76,     0,    89,    59,     0,    21,     0,   230,   106,     3,    74,   152,   205,    11,   205,   221,   222,   169,   161,    59,    99,   111,     0,     1,    26,   193,     6,   158,     4,   235,   203,     0,   121,    83,    75,    61,    52,   217,     0,   196,   103,   245,    87,   214,   247,   175,   141,     0,   207,   229,    66,    61,   160,   156,   249,     3,   130,   187,   245,    84,   130,    20,   208,    24,   238,   128,    47,    42,    87,     0,   105,   104,   236,     0,    55,    95,    69,   249,     0,   122,   107),
   (    8,    17,   145,   209,    80,   184,    23,   132,     0,     0,    33,   129,   245,   183,   177,    37,   114,   115,     7,    18,   190,     0,   141,   219,    34,    10,   172,     0,   245,   229,   119,   191,   145,   159,   104,     0,   114,   243,   221,   143,    66,     0,   251,   157,   108,   143,     2,   178,    23,   209,   166,   123,    43,   124,   247,    86,     0,   244,    55,    49,   119,     0,    54,    24,    60,   162,    44,   239,   175,   166,   246,     0,     0,   226,   148,   172,   105,    16,   104,    61,    27,    51,   227,    40,   134,    43,    70,   224,   189,   248,   232,    39,    18,   124,    35,    57,   166,   176,    54,    53,     0,    98,   180,   245,     5,    18,   154,   169,   166,   202,     0,    65,    95,   147,     3,   112,   218,   222,     0,   160,     8,   145,    85,    36,     0,   119,   149,   213),
   (  171,    45,    99,    75,     5,    91,    62,    11,    95,   248,    85,    34,   133,    67,   152,    13,   220,   236,   193,   168,   146,   141,     0,   143,   252,   251,   197,   147,   191,   255,     0,   179,   192,   239,   219,    32,     0,   107,   159,   196,     0,    63,   223,   194,    63,    83,   166,    19,   235,   215,    17,    40,    48,     6,   140,   242,    43,   129,    45,    34,    67,    32,    52,   150,   236,    56,   168,    37,   188,    84,   114,    81,     0,   158,   103,   185,   184,   176,   105,   142,   138,   239,     8,   220,   161,    46,   159,    57,   245,   190,   109,    60,   173,    13,   242,   211,    18,   177,    59,    61,     0,   217,   114,    35,   223,   159,    66,   228,     0,    29,   107,    69,    24,   119,   225,   184,   111,   101,   121,   111,   175,   169,     0,   132,   205,     0,   101,   212),
   (    1,   126,   253,   116,    77,   133,   212,     0,   147,     0,   121,   195,   156,   252,    78,    60,    44,   134,   103,    97,   181,   219,   143,     0,   125,   241,    56,    63,   121,   128,     9,    24,    44,    35,    75,    50,   117,   169,    90,    91,   109,   149,    52,    93,   120,     2,    17,   108,    19,   202,   198,   186,   105,    86,   237,     0,    29,    90,   213,   167,    92,    51,     0,    32,   152,    98,   249,    48,   144,   119,    56,   253,   122,    59,   113,     0,    63,   230,   178,   167,   145,   229,   234,   152,   105,   252,   226,    46,   143,   174,    99,   227,   117,   196,   248,   148,    62,    76,    27,    89,     0,    91,   249,    27,   195,    59,    61,   235,   236,    31,     0,   145,   150,   158,    44,   148,    74,     0,   136,    73,   200,   142,   137,    83,   207,   158,     0,   216),
   (  213,   213,    23,     1,   253,   229,   114,    71,    62,    66,    15,    48,    66,    82,   183,   144,   115,   103,   108,     0,   130,    34,   252,   125,     0,   236,    28,   166,   142,     8,   181,     0,   160,    71,    13,   208,   153,    16,    56,   224,    52,    58,    43,   113,   105,    57,    59,     9,    27,     0,   201,   125,   171,   235,   211,   115,     0,    33,    44,    73,   205,   232,    98,   204,   142,   246,   206,    24,   243,    69,   136,   194,    37,   255,   229,   208,     0,   212,    77,    85,   124,    96,    86,    53,    93,   253,    72,   149,   243,   111,   155,     0,   103,    69,   171,   227,   177,   110,     8,     0,   207,    67,   227,   165,    21,    58,    54,   166,    31,    16,    22,    13,   129,    33,    27,   139,    33,   132,    22,   215,   107,     0,     5,    85,   210,   107,    99,   252),
   (    0,    60,   208,   103,   197,    88,   100,    79,   100,    73,   139,   215,   109,   158,   118,   140,   118,    91,   196,    97,   213,    10,   251,   241,   236,     0,    68,    18,   209,    89,   198,   195,     0,   128,   105,   186,   179,   185,   123,   112,     0,   240,   250,    79,   253,   151,   160,    63,   147,   175,   184,   234,    42,   226,    26,    16,    30,    54,   180,     0,    72,    16,    94,   160,    35,   153,   234,     0,   157,    78,   243,    81,    62,   236,   180,   101,     6,     0,    16,    94,    59,   169,    16,    58,   236,   234,    29,   209,   120,    95,   207,   227,     0,   184,   174,    93,   128,   252,   150,   160,   138,    32,    20,   240,   193,   237,     0,   251,   254,   177,     0,     9,   194,   205,   255,   178,   212,    41,   231,   163,     0,   211,   125,   159,   199,    34,    74,   169),
   (  142,   217,   178,   110,    94,    52,    16,   108,   109,   166,    36,    93,    49,   239,    26,    83,   191,   215,    54,    98,   176,   172,   197,    56,    28,    68,     0,    80,   145,   176,    62,     0,   245,   239,    87,     0,    21,   151,   230,   193,   101,   194,    94,    79,   180,   174,   186,     6,   127,   212,    89,    67,     0,    81,    86,   124,     0,    92,   151,   232,   225,    25,   167,    63,    30,    80,    77,   231,    20,   160,   252,   243,   232,     0,   213,   182,   170,    22,   243,   100,   223,   128,     0,   254,   100,    48,     0,   102,    29,   238,   197,   235,   235,   146,   227,   241,   215,   154,   146,     0,    79,   100,     0,   217,    98,   148,   100,    42,     0,     0,   148,    46,   248,   231,   111,     0,   135,   214,     0,    38,   113,   233,     0,     0,   174,   174,   231,   231),
   (  131,     0,    18,    87,   220,   161,    28,     1,   251,   225,   144,     3,   154,   177,    87,   157,    64,   182,    39,     0,   253,     0,   147,    63,   166,    18,    80,     0,   107,   155,    35,   230,   121,     0,    73,    42,    43,   195,    55,   241,    64,   211,     2,   209,    96,   140,    70,     0,   123,   207,    73,    18,   240,     0,   182,   141,   191,   111,    10,     0,   144,    86,   235,   119,   166,   140,   209,   203,    95,     5,    60,    41,   187,   148,   241,   212,   119,    69,   193,   163,   165,   135,    32,    53,   132,     0,     0,   142,   235,   170,   195,    20,    93,    16,     0,   199,     0,   211,    91,     6,   151,    59,   131,   240,    34,   211,   223,     8,   164,   114,   139,   238,    16,   187,   203,    71,     0,   210,   124,   195,   239,   240,    97,    14,    59,   113,   244,     0),
   (    0,   203,    99,   141,    57,   191,   190,   204,   255,    79,   133,   135,    66,   119,   158,   219,   115,     0,   135,    95,   216,   245,   191,   121,   142,   209,   145,   107,     0,    77,   147,    32,   216,     0,     7,   249,    28,   251,   179,    83,   186,   221,   218,    43,    67,   105,   233,     0,   249,   237,   196,   179,    61,   100,   130,   218,   154,   243,    75,   178,    71,   240,   185,   226,   159,   138,     0,    42,   174,   246,   152,   233,     0,   197,   242,    47,    40,   137,    10,   136,    24,   236,   205,   169,   138,    63,     0,   192,    12,    53,   157,     0,    33,    29,    35,   196,   251,   139,   113,   144,   150,   254,    16,   146,    82,   183,    77,   252,    81,    74,   136,     1,    29,   105,    77,     0,   192,   115,   104,   191,   225,     0,    20,   243,     0,    52,     5,     0),
   (  184,    55,   166,   201,   156,     0,    39,   136,    47,   152,     0,   201,   100,    74,    96,   210,    63,   191,     0,    70,   218,   229,   255,   128,     8,    89,   176,   155,    77,     0,    41,   103,   138,   132,    33,   248,    57,    73,    85,   211,   151,    84,   145,   214,     0,    32,   103,   240,    92,   123,   154,    27,    35,   170,     0,    83,    58,   219,     5,   220,   110,    25,     0,    71,   157,   211,   251,    80,   194,    11,   133,    12,   161,    71,    44,   157,   152,    97,    52,   180,    94,   149,   161,    30,     4,   153,   244,   202,   101,   215,   186,   195,    39,   230,   134,    43,     0,    29,     0,   179,   254,   190,     0,   238,    84,   232,     0,    71,   239,   203,   162,   133,    93,    25,   217,    62,    70,     7,    53,     0,   162,     3,    55,    74,    12,    27,     0,    99),
   (   80,   125,   202,   239,    61,   162,   145,   145,    21,   233,   135,   167,   231,   188,    24,   112,   201,    82,   123,    66,   234,   119,     0,     9,   181,   198,    62,    35,   147,    41,     0,    28,   109,   170,    16,    51,   119,     0,    41,     0,   149,     0,   165,    97,     1,     0,   105,   186,   233,   151,    14,     1,    54,     0,     0,   136,   134,   184,    31,   123,   115,   115,   154,   237,    28,   134,   169,   141,   221,   191,   249,    85,   124,    61,   238,   156,   107,   153,   134,     7,    83,    96,   137,    77,   158,    26,   225,   113,   199,   126,   170,    95,   181,   239,   123,   153,    61,     0,   102,    36,     0,   239,   158,    22,   160,   116,   249,   217,   214,   254,   200,   197,   106,    93,    78,     0,   196,   144,     0,    70,   139,    77,     9,   136,   117,    39,    72,   165),
   (   98,   202,   248,    81,    39,   159,   218,     5,   232,     0,     0,    71,    47,   158,    39,   168,   100,    11,   162,   181,   153,   191,   179,    24,     0,   195,     0,   230,    32,   103,    28,     0,   162,   229,   129,   178,    94,    31,    29,     6,    99,     0,    28,    47,   126,   174,   209,   206,   234,    48,    14,    62,     0,   160,     0,   149,    44,   138,    72,    28,   167,    70,    68,   195,   204,   235,   100,   218,    71,    56,    32,     4,   232,     7,    50,    88,   129,    24,   192,    76,    68,    10,    37,   108,   219,     0,   250,   151,   139,   204,   241,   186,   100,    83,    89,     0,   253,   233,   228,    26,   145,    61,    33,   180,   228,   167,   146,     0,   188,    84,    37,   191,    37,     2,   249,    67,    61,   224,   103,   100,   102,   119,   115,    43,   117,   178,     0,   191),
   (  124,   209,     2,   246,    60,   242,    69,   232,   250,    92,   208,     1,   141,   139,   204,    62,   145,   213,    77,   104,   252,   145,   192,    44,   160,     0,   245,   121,   216,   138,   109,   162,     0,    14,    12,     0,     0,   255,    27,   247,   234,    34,     0,     0,   146,   162,     9,   217,     4,    64,   192,    34,   207,   170,    13,    19,   142,    40,   136,   107,    84,    57,    19,    24,   227,   207,   116,     0,   253,   150,   238,   253,     2,   171,   249,   119,   235,    75,   226,   144,    63,     0,   138,   164,   204,   138,   243,   198,   195,    88,    45,   108,    45,   191,   168,   209,   100,   214,    82,   203,     8,     0,   108,   116,   160,    87,   127,   125,    91,   172,   144,   198,   197,     0,    17,   140,    25,   249,   211,    64,   191,   208,   197,    28,    23,    72,   246,   245),
   (  139,   251,   170,     0,    37,     0,    60,    19,     0,    66,    28,   156,    21,     0,    83,    47,   102,   192,   180,     6,   120,   159,   239,    35,    71,   128,   239,     0,     0,   132,   170,   229,    14,     0,   163,     7,    83,   172,    56,   159,     0,   245,   155,   212,   124,     0,   174,   187,    70,   178,   213,    91,   205,   146,   154,   203,   109,    26,   106,    87,   216,     3,   163,     6,    56,    93,    67,   177,   229,   213,     0,    17,    80,   107,   176,   222,   245,    67,   243,    70,   127,    30,   180,    11,   170,   103,   211,    73,     0,   191,   249,   112,   170,    60,     0,   167,     8,     0,   233,   135,   171,   101,    93,   139,   121,   159,   129,   104,   204,    31,     0,   153,   238,   211,    41,   175,     0,   230,   113,   106,    60,   201,   104,   155,   117,    39,   176,     0),
   (  146,    48,    59,   230,   248,    66,   183,    31,    22,     0,   117,   184,    40,    76,     0,   211,   103,    25,    56,    95,   202,   104,   219,    75,    13,   105,    87,    73,     7,    33,    16,   129,    12,   163,     0,    52,   152,    77,   187,     0,   173,   179,   181,   128,   245,   168,    45,   137,     7,   253,     0,    11,   131,   176,   187,    86,   230,    16,   138,     0,    97,   188,   210,   138,   142,   183,     0,   105,     3,    98,     4,   109,   252,    77,    85,    31,   205,    44,   131,   194,   104,   149,   248,   125,   137,    72,     0,   147,   173,   211,   211,     0,   229,   191,    76,   207,   146,    13,   123,   207,   238,   227,   222,   129,    80,    61,     7,   210,    51,    32,    28,   244,     0,   164,   104,    96,    64,   205,    86,     0,    20,     0,    74,   139,   152,   157,    57,   151),
   (   47,   171,   140,   119,   183,    64,     0,    55,   137,    48,    70,   153,     9,    91,   123,   185,   194,   141,    19,   242,   161,     0,    32,    50,   208,   186,     0,    42,   249,   248,    51,   178,     0,     7,    52,     0,     0,     0,   116,   235,    32,     0,    38,    74,   114,   133,   153,    16,   134,   119,    46,     0,   184,   219,   105,    46,     8,    47,   113,     4,     2,    96,   228,   244,     0,    53,   177,   158,    48,    47,    55,   254,    33,   250,   154,   113,   168,    83,   118,   170,     0,    91,    78,   253,     7,   127,     8,     0,   109,   183,    70,   158,    43,   104,   183,   158,    82,    12,   141,    98,    68,   154,     0,   232,    42,   141,     0,   234,    75,    68,    68,     0,    46,   173,   237,   236,   251,     0,     0,    81,   131,   238,   231,   193,   234,   119,    79,    96),
   (  220,    95,   220,   166,    15,    63,    60,    42,   171,     0,   110,   189,    13,   211,   156,   244,   166,   221,   148,   106,   245,   114,     0,   117,   153,   179,    21,    43,    28,    57,   119,    94,     0,    83,   152,     0,     0,   121,    65,   109,   181,    61,    28,     2,   215,   178,    73,   255,    26,   181,   246,   241,    39,    34,   226,   209,   132,   202,   199,   157,   249,   225,   241,   144,   200,   235,   198,    67,   197,   210,   196,    65,    50,   124,   176,     0,    62,    58,    23,   109,   207,   166,   116,   144,   206,   187,   163,   247,   148,   166,   200,   156,    31,   180,     8,   142,   149,   106,   228,    56,    80,     0,    34,     9,     4,    84,    98,   211,    46,    81,   253,   244,    56,     1,   203,   100,    32,     0,     0,   219,   110,   154,   167,   248,   254,    98,   152,     6),
   (    0,    57,   212,     0,    86,   213,   211,   137,    51,   142,   247,    70,   225,   173,    24,   231,     0,   200,    14,   129,    78,   243,   107,   169,    16,   185,   151,   195,   251,    73,     0,    31,   255,   172,    77,     0,   121,     0,   154,   116,    21,     2,   245,   211,    42,    23,   106,    75,    43,     8,   171,    38,   110,    64,    80,    67,    91,   159,     0,   197,    72,    23,   191,    60,    40,   199,     0,   249,    41,   151,    37,   119,    96,     5,   122,     3,    60,    12,   159,   233,    82,   140,   115,   232,   103,   185,    19,    27,    81,     0,   251,    36,    36,     0,    15,   148,   141,   134,     0,   206,   209,   192,   141,   237,   247,   131,   109,   250,    65,   224,   140,   174,    88,   120,   214,    75,   145,   139,   143,     0,    95,   248,   168,    19,   205,   181,    98,   219),
   (  129,   101,    93,    75,   117,   218,     0,     0,   122,    24,    81,    54,   116,   240,    90,   130,   202,   155,    82,     0,    81,   221,   159,    90,    56,   123,   230,    55,   179,    85,    41,    29,    27,    56,   187,   116,    65,   154,     0,   159,    26,   238,     0,   248,    94,    38,    73,    68,    13,    29,    78,   235,   232,   188,   175,   186,    17,   165,   235,     0,   211,    31,   248,    75,   127,   230,   198,   231,    70,   156,   201,   132,   197,   255,   218,   221,    33,   199,   139,   129,   230,     7,    50,   199,    12,   178,   121,   152,    38,   110,   252,    37,   213,    22,   126,   140,   236,     3,    72,   221,   135,   198,    33,   115,   122,   234,   255,   238,   148,   103,   135,     5,   239,   174,    65,    76,    74,   130,    45,   157,    62,    29,    74,    86,     0,   246,   169,   169),
   (  198,   214,     3,   204,    68,   147,    98,    80,    66,     0,    94,   199,    93,    13,   234,    66,   226,   237,    78,    19,    65,   143,   196,    91,   224,   112,   193,   241,    83,   211,     0,     6,   247,   159,     0,   235,   109,   116,   159,     0,   148,   117,     0,   204,     0,   116,   130,    19,   124,     0,   224,    29,    25,   147,   191,    50,     0,   225,   203,   205,    92,   149,   250,   114,   160,   172,   226,     0,    31,    72,   153,   232,    94,   236,    60,   133,    45,   166,   236,   151,   180,   141,     1,    28,    59,    82,    57,   134,   253,    32,   231,   144,   158,   165,    36,     0,    81,   167,   208,   204,    24,   118,   228,   127,     0,   131,   123,   175,    53,     0,   237,   120,   222,   113,    27,   164,   226,    91,    98,    71,   181,    24,   137,    89,   203,   138,    51,    86),
   (   63,   155,    77,    25,   207,   198,   197,    75,   142,   219,   191,     0,   145,    70,   209,   151,   198,   222,    59,    26,   225,    66,     0,   109,    52,     0,   101,    64,   186,   151,   149,    99,   234,     0,   173,    32,   181,    21,    26,   148,     0,    10,   222,    69,   165,   213,    47,   189,   140,     0,    72,     0,   145,   129,     0,    51,     0,    33,    53,   204,   114,    64,    21,    79,    22,    63,   182,    88,   152,   120,    24,   191,   162,   171,   253,   137,    77,     0,    29,   231,   245,    38,   178,     8,   148,   218,    58,     1,     0,     0,   207,   140,    62,     0,   133,   235,   126,   180,   225,   214,   169,   220,     0,   101,   195,    18,    56,     0,    43,   171,   220,   153,    51,   200,    43,   115,    93,    80,    35,    60,     0,   159,   167,   107,    54,     0,   143,   236),
   (   36,    57,   142,   213,    77,   105,   108,   202,    52,   135,   252,   202,   155,   182,     0,   168,     0,   152,   101,    71,   212,     0,    63,   149,    58,   240,   194,   211,   221,    84,     0,     0,    34,   245,   179,     0,    61,     2,   238,   117,    10,     0,     0,    55,   180,     1,   115,   140,   185,   250,   234,   200,   106,   108,     0,    30,   216,    64,   237,   246,   147,   202,    28,    40,     0,     0,   101,   176,    59,    32,   185,   190,   128,   136,   221,   179,   193,   201,    19,     0,   185,   164,   214,     2,    61,   139,   230,   156,   125,   195,   239,   118,    89,    30,   132,   195,    69,   218,    36,   209,    37,   203,   255,    50,     0,   128,   176,   211,   192,    39,    66,     0,   217,   223,   238,    27,   180,    76,   193,     0,     2,   149,   130,   141,    13,   194,   152,    28),
   (  117,    82,    46,    78,    25,    44,   132,     0,    82,   240,   233,   105,   247,   195,    93,     0,   101,     0,    10,    22,    86,   251,   223,    52,    43,   250,    94,     2,   218,   145,   165,    28,     0,   155,   181,    38,    28,   245,     0,     0,   222,     0,     0,    88,   147,   208,   239,    88,    52,     0,   221,   158,    92,    75,   110,     9,    24,   148,     0,   119,    49,    74,    53,    25,   245,   213,    74,   188,   118,    83,   118,    33,     0,   123,   216,    91,   209,    35,   111,   220,     0,    52,   137,    34,    18,     3,   118,   148,    53,   199,   145,   178,   149,   124,   213,    96,   233,   110,   193,    31,   148,    29,    78,   185,    37,   219,   105,   178,   169,   234,     0,   203,   128,    53,   147,    28,     0,   150,     2,   155,   197,   134,   176,    48,   200,    98,   221,    27),
   (  219,   173,   186,    75,    71,    17,     9,   206,   186,   214,   148,    25,   214,     0,   104,   149,    82,   223,     0,   182,     0,   157,   194,    93,   113,    79,    79,   209,    43,   214,    97,    47,     0,   212,   128,    74,     2,   211,   248,   204,    69,    55,    88,     0,   139,    63,   143,   170,   133,   160,   149,   178,   110,    30,   122,   223,     9,    57,   100,   124,   254,    72,   182,   143,    74,   157,    13,   158,     0,   202,   178,   202,     0,   233,   237,   172,   159,    77,    67,    34,   150,   197,    72,   140,    57,   255,   207,    15,   237,   202,   205,     0,    78,   241,   210,   185,   152,   115,   117,   121,   199,   106,    68,   149,    46,   113,    14,   248,    55,     0,     0,    99,   225,    47,   156,   127,   239,   112,    19,   231,    69,    88,   152,    46,     0,     0,   218,   148),
   (   38,   169,     0,   122,   109,   204,   147,   193,   132,   219,   159,   206,     8,    98,    22,   200,    51,   120,   186,    72,   152,   108,    63,   120,   105,   253,   180,    96,    67,     0,     1,   126,   146,   124,   245,   114,   215,    42,    94,     0,   165,   180,   147,   139,     0,    54,    68,   153,   229,   133,   236,   238,    84,     0,     0,   188,   214,    51,    14,    43,     0,   123,    79,     7,     3,    32,    78,   168,   254,   212,   224,   122,     0,    69,   243,    70,    22,     0,    75,   198,   203,   146,   247,   127,    59,    63,   226,    24,     3,   109,   207,   223,   100,     0,     0,   116,   113,   210,    61,   108,   189,    74,   221,   124,    74,   199,    46,    67,    83,     0,   228,    88,   250,   201,     6,   109,   242,   141,   139,   103,   237,   235,     0,    94,    25,     0,     8,    23),
   (  198,     0,   230,    68,     0,    64,     0,   253,   201,   107,     0,    89,   158,   121,    47,   210,   183,   193,   210,    15,   231,   143,    83,     2,    57,   151,   174,   140,   105,    32,     0,   174,   162,     0,   168,   133,   178,    23,    38,   116,   213,     1,   208,    63,    54,     0,   223,    46,   127,   189,   100,     0,    37,     0,   189,    70,   118,     0,    41,   122,   121,    14,   182,    53,   116,   158,   172,    96,    20,    43,   219,   202,   118,   121,   196,     0,   177,   131,    16,   238,    31,   253,    26,   184,    69,   190,    19,   244,   174,   217,    97,    93,   186,   106,   139,    80,     0,   230,   237,   177,   198,   212,   121,   206,   109,    14,   250,     0,    44,    47,   151,     0,    41,     4,   127,   168,    84,     0,    60,    79,   197,   230,   156,   210,    83,   165,    42,   133),
   (  212,   170,    24,    38,   146,   114,   166,   169,   223,   103,   107,    57,     0,     5,   246,   184,    79,   210,    96,    37,   123,     2,   166,    17,    59,   160,   186,    70,   233,   103,   105,   209,     9,   174,    45,   153,    73,   106,    73,   130,    47,   115,   239,   143,    68,   223,     0,   137,   219,   177,    19,   222,   248,   130,   161,     0,   254,    96,     0,   237,   221,    15,   207,    85,   241,   210,   182,     0,   152,   211,   137,   116,   122,    12,   163,   247,   221,    73,    96,    42,    41,   229,    39,   132,    42,    36,    33,   102,    57,    67,     0,   143,   246,    29,   234,   115,    76,   114,     0,    63,   229,   254,   222,    78,    96,   245,   236,     0,    49,   168,    74,   171,   210,   167,    51,    27,   220,   138,   132,    24,     0,   112,   151,   218,   146,   215,   135,   253),
   (  184,    64,    48,     0,   149,   211,     5,    11,    91,   217,    34,     0,    90,   117,   189,   178,    18,    44,     0,    83,    76,   178,    19,   108,     9,    63,     6,     0,     0,   240,   186,   206,   217,   187,   137,    16,   255,    75,    68,    19,   189,   140,    88,   170,   153,    46,   137,     0,    30,   153,   228,   188,   152,   234,   253,   158,   172,    19,    74,    71,   150,    33,   176,    33,   145,     5,     1,   174,   176,   222,     0,   139,   176,   158,   163,    72,   146,     9,     0,   185,     0,   219,    38,   238,    71,   231,   100,   164,     0,   236,   196,    52,     1,   244,   190,   198,   135,    61,    88,   170,   130,     0,   116,   233,    50,   196,   120,    32,   178,    97,   169,    92,     0,   132,    44,   152,   184,   236,    40,   167,    72,   145,    37,   134,   252,   140,   117,     0),
   (   29,    42,   232,    33,    25,    69,    81,    30,     0,   252,    15,   130,    50,   134,   236,    94,   162,     0,     0,    24,     0,    23,   235,    19,    27,   147,   127,   123,   249,    92,   233,   234,     4,    70,     7,   134,    26,    43,    13,   124,   140,   185,    52,   133,   229,   127,   219,    30,     0,    16,   206,   255,    20,     0,    77,     0,   185,   224,   252,    82,   121,   137,   189,   193,   133,   145,   170,   244,    87,    98,   240,    10,   220,   121,   182,   160,    77,   112,    17,   141,   119,    24,     0,    52,   237,   207,   108,   201,    85,   133,   229,    24,    52,   234,    54,    80,   210,   197,    85,    51,   190,   168,     0,   116,    25,    46,   160,   223,     0,    40,   249,   253,    17,    11,    33,   253,   199,    96,   109,     2,   175,    13,     0,     5,    42,    80,   167,   243),
   (  123,   135,   205,   249,   210,    49,   230,   231,   201,   236,    67,   152,   162,   159,   149,   141,   137,    94,     0,    84,    89,   209,   215,   202,     0,   175,   212,   207,   237,   123,   151,    48,    64,   178,   253,   119,   181,     8,    29,     0,     0,   250,     0,   160,   133,   189,   177,   153,    16,     0,    67,    50,   188,   114,   128,   120,   246,   240,   169,   198,   163,   113,   206,   232,   224,   222,     0,   203,   145,     2,    24,    47,   186,    17,   118,    83,    61,    80,    82,   196,    90,   173,   130,    10,   191,   229,    86,   138,    32,   239,    68,   105,   214,   196,   116,   173,   161,   134,   182,    56,   123,   195,     0,     0,   163,    33,   224,   182,   125,    52,   165,   134,   112,   197,   137,     2,   112,   211,    29,    12,    59,   244,   200,   215,   206,    58,    51,    36),
   (  248,     0,    70,   231,   253,   137,    18,    70,   150,   159,   157,    25,    59,   143,   237,    83,    98,   112,   167,   137,    59,   166,    17,   198,   201,   184,    89,    73,   196,   154,    14,    14,   192,   213,     0,    46,   246,   171,    78,   224,    72,   234,   221,   149,   236,   100,    19,   228,   206,    67,     0,    42,   131,   199,    74,   173,   213,   158,   225,    46,     0,   162,   255,   206,    83,   232,     0,    32,    61,    71,    82,   216,   183,   133,   145,   219,   149,    99,   211,    58,   102,   205,   196,   167,     0,    47,    94,    51,    69,    52,   104,     0,   234,     0,    49,    51,   248,   191,   226,     0,     5,   161,    32,   177,   110,   124,   205,   162,   177,    26,   205,    31,    18,    68,    76,    11,    11,   144,    66,   130,    77,   165,   225,    22,   183,   136,     2,   237),
   (  192,    29,   239,    76,   102,   156,   184,     4,     0,    94,   149,     0,   190,    73,   224,   100,   157,    96,   168,     1,     0,   123,    40,   186,   125,   234,    67,    18,   179,    27,     1,    62,    34,    91,    11,     0,   241,    38,   235,    29,     0,   200,   158,   178,   238,     0,   222,   188,   255,    50,    42,     0,   239,   214,    43,    44,   239,   206,     0,    18,   133,    40,    48,    67,   220,   174,    75,    17,    32,    73,    13,   154,   186,    41,   235,   214,    67,   143,   233,     0,    77,   237,    68,    44,   135,   183,    49,    84,   164,   142,   145,     0,    20,    39,    80,    18,   244,    61,   238,    96,    87,   164,     0,    71,   194,    19,    62,   173,    10,   236,    78,    29,   140,    49,   159,    49,   131,    71,   150,   124,   239,   223,    29,    30,     0,   106,     1,    24),
   (  224,   234,   118,   157,     4,   236,    55,     0,   236,   146,     0,   181,   129,    69,     0,   209,    80,   197,   187,    21,    21,    43,    48,   105,   171,    42,     0,   240,    61,    35,    54,     0,   207,   205,   131,   184,    39,   110,   232,    25,   145,   106,    92,   110,    84,    37,   248,   152,    20,   188,   131,   239,     0,   228,    22,     0,   199,   179,    67,     0,    31,    56,   250,   199,   225,    24,   253,   158,   184,     0,   139,   235,   116,   207,   127,     0,    73,   181,     0,   162,   216,   191,    83,     6,     9,   235,   169,    23,    58,   244,    67,   235,    63,   148,   189,   205,   253,    54,    86,   168,    33,   211,   223,   144,     0,     0,   217,    73,   141,     0,    11,     0,   209,   210,   154,   149,   183,   166,    41,   230,   222,     9,   199,   193,   131,     0,    81,     0),
   (  172,    83,    29,    41,   110,   181,   199,    51,   252,    44,    43,   111,    73,    61,    32,   155,    63,   157,     1,   131,     0,   124,     6,    86,   235,   226,    81,     0,   100,   170,     0,   160,   170,   146,   176,   219,    34,    64,   188,   147,   129,   108,    75,    30,     0,     0,   130,   234,     0,   114,   199,   214,   228,     0,    35,   119,    40,    80,   128,    20,    60,   113,   227,     0,     0,    99,   129,   237,    20,   230,   110,   146,     4,   243,   233,   198,   225,    74,     0,    12,   131,   253,   225,   125,    55,    87,     0,   200,   211,    31,    33,   100,   141,   241,   185,   203,   252,    84,   109,   246,    78,    37,   242,   202,     0,   128,   187,   138,     0,    48,     0,    35,    65,   240,   205,   106,     1,    83,     7,    61,    13,    19,   133,   222,   218,   153,    13,   169),
   (    7,   165,   140,   204,   233,     0,   131,     2,   179,   169,   245,   252,   137,    25,   111,   100,    92,    27,    65,   179,   230,   247,   140,   237,   211,    26,    86,   182,   130,     0,     0,     0,    13,   154,   187,   105,   226,    80,   175,   191,     0,     0,   110,   122,     0,   189,   161,   253,    77,   128,    74,    43,    22,    35,     0,     0,   108,   199,    75,   234,     0,     0,   110,   236,    11,    23,   162,    59,   123,    64,   225,     0,    54,   115,   120,   218,     7,   149,   114,     0,   123,   206,     8,   164,    72,   113,    23,   206,    45,   237,   158,   113,    73,     0,   241,    93,    15,   164,   225,    25,    34,     0,    18,   218,    59,    23,   253,   194,    97,     1,   228,   132,   211,    38,   215,    69,     0,    14,   188,   107,    94,    94,    26,   110,   149,    67,    85,   196),
   (  130,   127,   175,   214,     1,   161,   167,   129,   216,    25,     0,     0,    88,   162,   254,    48,   168,   177,   206,    67,   106,    86,   242,     0,   115,    16,   124,   141,   218,    83,   136,   149,    19,   203,    86,    46,   209,    67,   186,    50,    51,    30,     9,   223,   188,    70,     0,   158,     0,   120,   173,    44,     0,   119,     0,     0,   202,     0,   114,   216,     0,   102,   217,    60,    24,    44,     0,   103,   150,   228,    85,    75,   223,    56,   131,    56,    27,    72,    17,     0,   194,   145,   102,    10,   237,    55,   148,   238,   103,    64,    34,   143,   203,   236,     8,   200,   135,   141,   220,   211,   242,   228,     0,   206,   210,   155,   139,   145,   103,    85,   243,   216,   175,   113,    46,    19,    38,   245,     0,   111,    89,   180,    59,   218,   105,    15,    15,    63),
   (    7,   237,   165,   213,    68,    30,   183,   235,   163,    48,   131,    74,    60,   130,   228,   110,     0,    52,     0,   166,     3,     0,    43,    29,     0,    30,     0,   191,   154,    58,   134,    44,   142,   109,   230,     8,   132,    91,    17,     0,     0,   216,    24,     9,   214,   118,   254,   172,   185,   246,   213,   239,   199,    40,   108,   202,     0,     0,   184,    39,   250,     0,   129,   154,   138,   191,   150,     0,    50,   215,   247,    88,    19,    50,   245,   194,   185,   212,   176,    77,    98,   182,   215,    28,   246,    79,   234,   100,    46,   188,    23,   162,     6,    20,   235,   137,   165,    41,   153,   255,   117,    46,    53,   220,   104,   234,   141,   111,    12,   182,     0,   149,   161,    73,   163,    30,   140,   230,     0,    30,   253,   153,   208,   216,   130,    89,    85,   222),
   (   68,    43,    43,   121,   181,     0,   143,    70,    57,    96,   195,   222,   107,    63,   152,    16,    52,   222,     5,   149,    74,   244,   129,    90,    33,    54,    92,   111,   243,   219,   184,   138,    40,    26,    16,    47,   202,   159,   165,   225,    33,    64,   148,    57,    51,     0,    96,    19,   224,   240,   158,   206,   179,    80,   199,     0,     0,     0,   193,   247,   134,    79,    30,    62,   184,     0,    75,    58,   180,    62,    49,    77,   249,   196,   208,   249,   115,    43,    90,   219,    63,    42,    36,   232,    17,   247,   114,     0,    46,    70,   254,   121,   255,     4,   247,   236,    64,    99,   157,   222,    69,   153,   219,     0,     0,   137,   181,   106,    49,   161,   149,   145,   163,   179,    21,   203,     0,   226,   146,   154,    29,   154,    96,   105,   116,   212,     1,   184),
   (   97,     0,   249,   141,   117,   172,   173,    39,   191,   109,     0,   159,   170,    23,   196,   184,   174,    34,    33,    58,   152,    55,    45,   213,    44,   180,   151,    10,    75,     5,    31,    72,   136,   106,   138,   113,   199,     0,   235,   203,    53,   237,     0,   100,    14,    41,     0,    74,   252,   169,   225,     0,    67,   128,    75,   114,   184,   193,     0,     0,   166,   233,     0,   173,   161,   213,   161,    17,    25,   241,   168,   178,   116,   229,   228,   182,     4,   227,    75,    62,    22,     0,    47,   232,   211,   118,    34,   253,    19,    77,   221,   214,    98,    86,   153,   150,    24,   248,    22,    32,    65,    54,    76,   205,   242,   102,    94,   250,   237,     0,    13,   242,    58,   215,     0,    26,   210,   181,    18,     0,   219,   194,     0,    47,    18,   187,    86,    16),
   (  198,    35,   196,    42,   168,   127,     0,    88,   134,   158,    43,   199,     0,   133,    60,   164,   102,   164,     0,   180,   205,    49,    34,   167,    73,     0,   232,     0,   178,   220,   123,    28,   107,    87,     0,     4,   157,   197,     0,   205,   204,   246,   119,   124,    43,   122,   237,    71,    82,   198,    46,    18,     0,    20,   234,   216,    39,   247,     0,     0,    85,    78,   241,   115,    28,    12,   254,   238,   119,    25,   125,   131,   150,     0,     0,   219,   137,   171,    87,    98,   128,   122,   188,   115,    83,   182,    28,   166,   245,    77,    80,    91,    61,   229,   238,    89,   168,   103,   252,   184,   233,   115,    12,   254,   124,    10,    20,   189,   230,    93,   218,   245,    98,   115,    33,    24,    79,   236,   152,   140,    40,     0,    93,    72,   110,   105,   185,   187),
   (   77,   113,   250,    75,    88,   184,   173,     0,     0,    95,   143,    92,     0,   118,   125,   187,   167,   180,    90,   235,    11,   119,    67,    92,   205,    72,   225,   144,    71,   110,   115,   167,    84,   216,    97,     2,   249,    72,   211,    92,   114,   147,    49,   254,     0,   121,   221,   150,   121,   163,     0,   133,    31,    60,     0,     0,   250,   134,   166,    85,     0,   156,     2,   151,    38,    13,   109,     0,    24,     3,   162,   148,   195,     0,    53,    96,   237,   107,   224,   255,    83,   231,   161,     0,   245,   184,   202,   227,   228,     7,    74,   214,     0,   122,   226,   156,   101,    70,   105,    35,   223,     0,    15,   241,    40,   201,   234,     0,   220,   199,   147,   155,   237,    39,   125,   232,    83,   182,   251,   227,   247,   164,   135,     0,   247,    64,    36,   101),
   (   49,   253,     4,    67,   164,    66,    33,   243,   223,    14,    62,   244,   163,   175,    96,   201,   160,    60,    10,    78,   205,     0,    32,    51,   232,    16,    25,    86,   240,    25,   115,    70,    57,     3,   188,    96,   225,    23,    31,   149,    64,   202,    74,    72,   123,    14,    15,    33,   137,   113,   162,    40,    56,   113,     0,   102,     0,    79,   233,    78,   156,     0,    25,   240,    52,   194,   237,    98,   125,    98,    22,     0,   232,   216,     9,   226,    96,   252,   189,   202,   192,   193,   206,   235,   185,   172,     0,     0,   145,   106,    66,     0,    59,    19,    92,   154,    50,    21,    25,   218,    96,   230,   235,   117,    23,   190,   178,   107,    43,   243,    89,     0,   181,   105,    30,     0,   230,    78,    48,   222,   208,   154,    92,    44,     7,    48,    25,     0),
   (  175,    48,    52,     0,   248,   125,   117,    97,   197,   196,    27,    50,    59,   115,    98,   129,    94,   124,   187,     0,   221,    54,    52,     0,    98,    94,   167,   235,   185,     0,   154,    68,    19,   163,   210,   228,   241,   191,   248,   250,    21,    28,    53,   182,    79,   182,   207,   176,   189,   206,   255,    48,   250,   227,   110,   217,   129,    30,     0,   241,     2,    25,     0,    34,    66,    77,   233,   232,   184,    28,     0,   203,   253,     0,    77,    79,     0,    28,   230,    16,    49,   144,    57,   159,     1,   140,   140,   122,    55,   127,   239,    73,    46,     0,     0,    29,   243,   156,    83,     0,   134,     0,    67,    73,   228,    55,    57,    95,    99,   242,   182,   176,    29,   214,     2,     0,   200,   143,   140,   120,    17,   178,   240,   158,   247,    30,   159,   196),
   (  202,    53,    73,   229,   129,    91,    15,     7,   186,    92,   157,   244,   104,   208,    93,   146,   221,    68,   250,    48,   222,    24,   150,    32,   204,   160,    63,   119,   226,    71,   237,   195,    24,     6,   138,   244,   144,    60,    75,   114,    79,    40,    25,   143,     7,    53,    85,    33,   193,   232,   206,    67,   199,     0,   236,    60,   154,    62,   173,   115,   151,   240,    34,     0,   115,   130,   231,   106,   238,   176,   176,    14,   199,    80,    47,   239,    58,    57,   141,   205,    79,   223,   185,   255,     0,     0,   210,    26,   220,   125,   120,   131,   244,    21,   233,   198,    77,   122,   205,   110,    88,   196,   112,    18,     0,   115,   195,    63,   174,   146,   129,   249,   113,   101,   163,   196,    55,    61,   146,     1,     0,   120,    99,   242,   161,   240,   240,   208),
   (    8,    53,   179,   183,   192,     0,    13,   153,   123,    77,   142,   145,    46,   204,    36,   233,   179,    11,   173,    27,   169,    60,   236,   152,   142,    35,    30,   166,   159,   157,    28,   204,   227,    56,   142,     0,   200,    40,   127,   160,    22,     0,   245,    74,     3,   116,   241,   145,   133,   224,    83,   220,   225,     0,    11,    24,   138,   184,   161,    28,    38,    52,    66,   115,     0,   209,    77,    38,   128,   217,   235,   252,   144,   125,   133,    98,    44,   205,   174,   148,   224,    22,   250,    93,     0,   147,    74,   226,   237,   153,   191,   125,     0,   227,   218,    49,   120,     0,    99,   223,    37,    45,    55,    88,   152,     0,   180,   161,    64,    81,   153,    32,     0,   125,     0,    63,   219,   132,   170,   130,    11,   101,   223,   133,     0,   119,    20,    83),
   (   39,     0,    63,    16,   175,    33,   248,   191,   133,    43,   255,    20,    97,    84,   239,    17,    41,    41,   254,    85,   161,   162,    56,    98,   246,   153,    80,   140,   138,   211,   134,   235,   207,    93,   183,    53,   235,   199,   230,   172,    63,     0,   213,   157,    32,   158,   210,     5,   145,   222,   232,   174,    24,    99,    23,    44,   191,     0,   213,    12,    13,   194,    77,   130,   209,     0,    15,    10,    21,    37,    63,     8,   121,   164,    54,    19,    71,    40,    51,    59,   161,   106,   205,   146,   245,   126,    90,   201,   131,   239,   238,     3,     0,   215,   131,   128,   162,   209,   126,     9,    63,   224,    58,     5,   210,     0,   249,    69,     6,    92,   103,    90,   186,    76,   237,   208,    94,   170,   107,    82,    52,    18,   254,   148,    23,    93,   227,   155),
   (  240,   239,   187,   157,   142,    72,   201,   101,   113,   178,    46,   153,   135,     0,    76,    50,    22,    78,    77,   126,    59,    44,   168,   249,   206,   234,    77,   209,     0,   251,   169,   100,   116,    67,     0,   177,   198,     0,   198,   226,   182,   101,    74,    13,    78,   172,   182,     1,   170,     0,     0,    75,   253,   129,   162,     0,   150,    75,   161,   254,   109,   237,   233,   231,    77,    15,     0,    87,    67,   130,   162,    62,    71,     0,    53,   155,    11,    92,    72,    80,   243,     0,     0,   192,   124,   252,   172,    79,    71,   145,    64,   220,   156,   202,    46,    12,   114,    85,    64,     0,   133,   127,   203,    62,   254,   134,   158,    27,   204,   185,   125,    24,   199,   181,   255,    98,   214,   223,    34,   203,   177,    38,   212,   115,    49,   165,   134,   250),
   (  185,     3,    18,   184,   122,    21,   168,    47,   157,   247,   248,     7,    95,   223,   159,    23,   230,   138,   122,    30,    99,   239,    37,    48,    24,     0,   231,   203,    42,    80,   141,   218,     0,   177,   105,   158,    67,   249,   231,     0,    88,   176,   188,   158,   168,    96,     0,   174,   244,   203,    32,    17,   158,   237,    59,   103,     0,    58,    17,   238,     0,    98,   232,   106,    38,    10,    87,     0,   238,   234,   127,   147,   201,   192,    90,    39,    85,   196,   179,   109,   152,     3,   183,   190,    79,    25,   125,     0,   188,   231,   248,    96,     0,    43,   186,    11,   137,   231,     0,    34,   201,     5,   146,    33,   172,     6,    21,    65,   132,     0,    92,    39,   191,   250,    50,   133,    82,   117,   111,    44,   211,    13,     0,     0,    33,   171,    22,    34),
   (  126,    64,    37,   113,    70,   250,    29,   219,    58,   123,   251,    26,     0,   251,   110,   235,    49,     2,     1,   173,   111,   175,   188,   144,   243,   157,    20,    95,   174,   194,   221,    71,   253,   229,     3,    48,   197,    41,    70,    31,   152,    59,   118,     0,   254,    20,   152,   176,    87,   145,    61,    32,   184,    20,   123,   150,    50,   180,    25,   119,    24,   125,   184,   238,   128,    21,    67,   238,     0,    35,   116,    30,   253,   183,   110,     0,     0,   168,    58,   153,   236,    78,     0,   246,   242,   246,   234,   247,   117,   191,   158,    56,    55,   105,   250,    78,   105,     0,   224,   178,   117,   248,   199,   208,   102,   236,   158,   125,     4,     0,    22,    20,    67,    92,    69,   207,   241,   194,    79,    38,   163,   228,   251,     0,    75,   230,   165,   181),
   (  131,    90,    36,   122,     0,   175,     0,     0,    65,   159,    61,   133,    87,    34,   203,    42,   112,    99,   165,   150,     0,   166,    84,   119,    69,    78,   160,     5,   246,    11,   191,    56,   150,   213,    98,    47,   210,   151,   156,    72,   120,    32,    83,   202,   212,    43,   211,   222,    98,     2,    71,    73,     0,   230,    64,   228,   215,    62,   241,    25,     3,    98,    28,   176,   217,    37,   130,   234,    35,     0,   158,     3,    80,     0,     0,    85,   233,    54,    40,   212,     1,   129,    15,   243,   169,    16,   142,     0,   211,    61,     7,   180,   213,   232,   160,   215,   162,   226,   149,    29,     7,   202,    81,   140,   133,     0,   168,    63,   203,   130,   153,   187,    91,    81,     7,   209,     0,     0,   204,     0,   241,    84,    12,   108,   225,   248,   243,     4),
   (   33,    40,     0,    80,   147,    79,     0,    57,    66,   172,   197,   177,   177,   186,   140,    94,   122,    86,   192,     2,     1,   246,   114,    56,   136,   243,   252,    60,   152,   133,   249,    32,   238,     0,     4,    55,   196,    37,   201,   153,    24,   185,   118,   178,   224,   219,   137,     0,   240,    24,    82,    13,   139,   110,   225,    85,   247,    49,   168,   125,   162,    22,     0,   176,   235,    63,   162,   127,   116,   158,     0,   188,   117,    17,   154,   199,   237,   181,    11,    16,   139,    27,   147,   149,    30,    68,    13,    42,   235,    23,   151,    41,   239,    57,    29,   152,   204,     9,     0,     0,    16,    98,    96,   187,     0,     0,   185,    58,   247,   203,   134,   176,   204,   244,   110,   177,    88,    14,   126,    55,   193,   171,    49,     0,   219,    67,   170,   107),
   (   62,    30,    82,   131,   161,   197,   131,   156,   232,   104,    25,    51,    85,   171,    37,   150,   113,   106,   238,    50,    26,     0,    81,   253,   194,    81,   243,    41,   233,    12,    85,     4,   253,    17,   109,   254,    65,   119,   132,   232,   191,   190,    33,   202,   122,   202,   116,   139,    10,    47,   216,   154,   235,   146,     0,    75,    88,    77,   178,   131,   148,     0,   203,    14,   252,     8,    62,   147,    30,     3,   188,     0,   128,     0,   183,    81,    72,   178,    56,     0,    23,   168,    55,    56,   121,   234,   139,   189,   253,   101,    34,    39,   224,    14,    52,   157,    58,   156,   148,    88,   161,     2,     0,    56,   245,   118,   197,    48,    52,   163,   193,   199,   140,    23,    36,    15,    36,   144,   174,     0,    34,   123,   183,    29,   112,     0,     0,    98),
   (  150,   244,    46,   177,   111,     0,    97,   106,   105,   160,   141,   152,    15,     0,    58,   141,    40,   102,   213,   110,   193,     0,     0,   122,    37,    62,   232,   187,     0,   161,   124,   232,     2,    80,   252,    33,    50,    96,   197,    94,   162,   128,     0,     0,     0,   118,   122,   176,   220,   186,   183,   186,   116,     4,    54,   223,    19,   249,   116,   150,   195,   232,   253,   199,   144,   121,    71,   201,   253,    80,   117,   128,     0,   186,    64,   198,     0,    97,     0,    24,     0,   230,     1,    65,   163,   143,   230,     0,   210,    17,   226,     0,    85,     0,   120,   108,     0,    51,   158,    14,    85,   232,     0,   119,    48,   207,    21,    35,    82,   216,   141,   192,   160,   147,    69,    35,   186,   179,   160,    85,   112,   192,   122,   248,   113,     0,     0,   157),
   (   96,    37,   136,     0,   146,   228,   193,   205,   104,     0,    18,   125,    52,   164,   108,   174,   119,   122,   175,   183,     6,   226,   158,    59,   255,   236,     0,   148,   197,    71,    61,     7,   171,   107,    77,   250,   124,     5,   255,   236,   171,   136,   123,   233,    69,   121,    12,   158,   121,    17,   133,    41,   207,   243,   115,    56,    50,   196,   229,     0,     0,   216,     0,    80,   125,   164,     0,   192,   183,     0,    17,     0,   186,     0,   106,   145,     0,   250,   156,   168,   131,   224,    92,   111,   123,    87,    87,    48,    17,   162,     0,     0,   110,   155,   239,    69,    51,    62,   116,     0,    13,    87,     0,   194,   175,   191,   253,   106,   169,   108,     0,   104,   206,   248,    87,     0,    49,   126,   209,   252,    69,   177,     7,    38,   204,   211,   251,     0),
   (  248,    24,   197,    62,   203,   250,    83,    54,   177,   162,   253,   135,   204,   110,     0,    79,     0,   179,   111,   110,   158,   148,   103,   113,   229,   180,   213,   241,   242,    44,   238,    50,   249,   176,    85,   154,   176,   122,   218,    60,   253,   221,   216,   237,   243,   196,   163,   163,   182,   118,   145,   235,   127,   233,   120,   131,   245,   208,   228,     0,    53,     9,    77,    47,   133,    54,    53,    90,   110,     0,   154,   183,    64,   106,     0,   128,   177,    71,   105,    23,   196,    14,   147,    80,   150,    40,    33,   241,   233,     0,    91,   187,    36,    50,   229,     9,   147,   199,   110,    11,     8,   100,   197,     0,   146,   246,   151,    55,   180,   171,    27,    27,   213,     0,   246,    20,    17,   228,   215,   161,   174,     0,    66,   233,   136,    68,   232,    41),
   (  102,   105,   124,   190,    51,   217,     5,    56,    70,   101,   142,     0,   155,   100,    62,     0,   158,     0,   241,   249,     4,   172,   185,     0,   208,   101,   182,   212,    47,   157,   156,    88,   119,   222,    31,   113,     0,     3,   221,   133,   137,   179,    91,   172,    70,     0,   247,    72,   160,    83,   219,   214,     0,   198,   218,    56,   194,   249,   182,   219,    96,   226,    79,   239,    98,    19,   155,    39,     0,    85,   199,    81,   198,   145,   128,     0,    60,   167,   175,   173,     0,   139,   137,    66,     0,     4,   183,   123,   232,    17,     0,   152,   173,   175,    47,   250,   199,    65,    89,     0,    65,   203,   120,    12,     8,    76,    55,   100,   243,   123,   146,   170,   246,   246,   208,   103,   152,     0,   116,    83,    96,   102,   104,     0,   181,   113,   180,   106),
   (  105,     0,   196,     3,   142,    51,   184,    76,     0,   188,    19,   201,   237,     0,   198,   214,   168,   233,     0,   173,   235,   105,   184,    63,     0,     6,   170,   119,    40,   152,   107,   129,   235,   245,   205,   168,    62,    60,    33,    45,    77,   193,   209,   159,    22,   177,   221,   146,    77,    61,   149,    67,    73,   225,     7,    27,   185,   115,     4,   137,   237,    96,     0,    58,    44,    71,    11,    85,     0,   233,   237,    72,     0,     0,   177,    60,     0,   144,     0,     0,   122,     0,   223,   120,   170,    65,   164,    57,    69,   122,    58,   109,     0,   106,   132,    58,   168,   204,   170,    71,    76,     7,   155,     0,    52,   129,     0,    10,     0,    83,   153,    24,   198,     0,   113,   219,    83,     2,   210,   131,    48,   196,     0,   217,   235,   154,   240,   122),
   (  245,   213,    89,    38,    46,   167,   247,   140,    47,    95,   121,   206,    63,   253,    52,   114,    25,    92,    39,    95,   203,    16,   176,   230,   212,     0,    22,    69,   137,    97,   153,    24,    75,    67,    44,    83,    58,    12,   199,   166,     0,   201,    35,    77,     0,   131,    73,     9,   112,    80,    99,   143,   181,    74,   149,    72,   212,    43,   227,   171,   107,   252,    28,    57,   205,    40,    92,   196,   168,    54,   181,   178,    97,   250,    71,   167,   144,     0,     0,    17,   183,   181,   255,   102,   244,   243,    64,   235,   211,    72,   148,     6,    97,   193,   156,    68,    22,    25,   216,    28,     0,    60,   176,   249,    29,   130,    27,   236,   102,   139,   141,    14,    43,   234,   191,   192,   175,    36,   253,   227,    56,   158,   190,   198,   250,   107,     3,   115),
   (   74,   200,   181,    63,     0,    95,    35,   215,   183,    23,    68,    68,   102,   192,   250,   234,   126,     0,   243,   227,     0,   104,   105,   178,    77,    16,   243,   193,    10,    52,   134,   192,   226,   243,   131,   118,    23,   159,   139,   236,    29,    19,   111,    67,    75,    16,    96,     0,    17,    82,   211,   233,     0,     0,   114,    17,   176,    90,    75,    87,   224,   189,   230,   141,   174,    51,    72,   179,    58,    40,    11,    56,     0,   156,   105,   175,     0,     0,     0,    92,    81,   175,   230,     0,     0,   126,   176,   114,    71,   190,    62,   239,    35,   112,    16,   129,   122,   131,    58,   252,    84,   181,   198,   159,    13,   187,   163,    94,   187,   156,    14,    39,   127,    99,    39,    86,   121,   198,    12,    27,     0,    29,    40,     0,   167,     0,   121,   250),
   (   25,   182,     0,   147,     0,    18,   183,   182,    10,     0,   176,   132,    72,     2,    25,   136,    91,    22,     0,    63,   121,    61,   142,   167,    85,    94,   100,   163,   136,   180,     7,    76,   144,    70,   194,   170,   109,   233,   129,   151,   231,     0,   220,    34,   198,   238,    42,   185,   141,   196,    58,     0,   162,    12,     0,     0,    77,   219,    62,    98,   255,   202,    16,   205,   148,    59,    80,   109,   153,   212,    16,     0,    24,   168,    23,   173,     0,    17,    92,     0,    54,   224,    58,    49,    83,   144,   212,   131,   107,   141,    72,    88,   252,   228,   163,   118,   139,    46,   238,    69,   229,   158,   186,   157,   191,    73,   251,    12,    17,    48,   133,     3,    60,   149,    86,    63,   118,     0,    90,   245,     0,    12,   145,   138,   151,    64,    84,   206),
   (  138,   103,    75,     0,    19,   226,   233,   155,   139,   113,    15,    64,   176,    94,    31,    93,     0,     5,   252,    32,    83,    27,   138,   145,   124,    59,   223,   165,    24,    94,    83,    68,    63,   127,   104,     0,   207,    82,   230,   180,   245,   185,     0,   150,   203,    31,    41,     0,   119,    90,   102,    77,   216,   131,   123,   194,    98,    63,    22,   128,    83,   192,    49,    79,   224,   161,   243,   152,   236,     1,   139,    23,     0,   131,   196,     0,   122,   183,    81,    54,     0,    99,   228,     0,     0,    91,    36,    46,    80,     0,   254,   210,   122,    61,   103,   224,   238,     0,     0,   253,   180,   248,   159,   154,    14,    95,   180,   140,   131,   178,    28,   142,   122,    53,    12,    21,   161,   254,   242,     0,   117,    61,   119,    34,    63,    66,    75,   163),
   (   55,   234,   178,   125,   240,    28,   134,   105,     0,   241,     3,   204,   140,   176,    71,    30,   212,   127,    48,   195,    75,    51,   239,   229,    96,   169,   128,   135,   236,   149,    96,    10,     0,    30,   149,    91,   166,   140,     7,   141,    38,   164,    52,   197,   146,   253,   229,   219,    24,   173,   205,   237,   191,   253,   206,   145,   182,    42,     0,   122,   231,   193,   144,   223,    22,   106,     0,     3,    78,   129,    27,   168,   230,   224,    14,   139,     0,   181,   175,   224,    99,     0,     0,   100,   140,   175,   162,   131,   253,    90,   233,   176,   166,     0,   192,   221,   187,   143,    97,    27,     0,   236,    48,   238,    64,   227,   100,   122,   187,   133,     2,    86,    51,    68,    37,     0,     0,    85,    13,     0,   157,    63,     9,    16,    13,   234,   132,     4),
   (   27,     0,    14,   199,   238,   117,   132,   251,    57,   231,    76,   162,   227,     0,     0,    59,   174,   153,   165,   211,    61,   227,     8,   234,    86,    16,     0,    32,   205,   161,   137,    37,   138,   180,   248,    78,   116,   115,    50,     1,   178,   214,   137,    72,   247,    26,    39,    38,     0,   130,   196,    68,    83,   225,     8,   102,   215,    36,    47,   188,   161,   206,    57,   185,   250,   205,     0,   183,     0,    15,   147,    55,     1,    92,   147,   137,   223,   255,   230,    58,   228,     0,     0,   228,   179,     0,    52,    37,    82,   244,   187,   139,   124,   115,   246,   139,   140,    34,   254,     0,    93,     0,   121,     0,     7,   134,    88,    19,   106,    90,   108,   114,    53,   201,   168,   224,   126,     0,   135,   100,     0,    55,    38,     0,   172,   188,   239,   246),
   (  160,   232,   216,   182,   104,    15,     0,   105,   137,   128,     0,   143,    53,   114,   228,   206,    47,     0,    62,   124,    52,    40,   220,   152,    53,    58,   254,    53,   169,    30,    77,   108,   164,    11,   125,   253,   144,   232,   199,    28,     8,     2,    34,   140,   127,   184,   132,   238,    52,    10,   167,    44,     6,   125,   164,    10,    28,   232,   232,   115,     0,   235,   159,   255,    93,   146,   192,   190,   246,   243,   149,    56,    65,   111,    80,    66,   120,   102,     0,    49,     0,   100,   228,     0,    72,    88,   229,   177,   200,    32,    70,     0,   103,    34,   193,   200,     0,   218,    68,    91,     0,    92,   240,     0,   177,    79,   175,   196,     0,   147,     0,   192,   247,     0,   255,    27,   238,   110,   195,   239,   128,    31,   247,   145,   130,    91,   210,    52),
   (   11,   214,   244,   107,     0,     0,    80,    30,   155,    27,    91,   178,     0,    56,   134,    46,    65,   105,    53,    65,   217,   134,   161,   105,    93,   236,   100,   132,   138,     4,   158,   219,   204,   170,   137,     7,   206,   103,    12,    59,   148,    61,    18,    57,    59,    69,    42,    71,   237,   191,     0,   135,     9,    55,    72,   237,   246,    17,   211,    83,   245,   185,     1,     0,     0,   245,   124,    79,   242,   169,    30,   121,   163,   123,   150,     0,   170,   244,     0,    83,     0,   140,   179,    72,     0,    71,   227,   211,    97,   154,     0,   248,   224,   194,     0,    36,   154,   160,    68,    55,     0,   114,   173,   171,   190,   206,    45,   129,     0,   201,   192,   125,    70,     0,   103,    85,   145,   168,    92,   124,    82,     0,   108,    39,   162,   245,   177,     0),
   (  128,    43,    83,   241,   194,   196,     2,   112,   150,   253,   114,   111,   151,   225,    33,   232,   254,   254,     0,    62,     0,    43,    46,   252,   253,   234,    48,     0,    63,   153,    26,     0,   138,   103,    72,   127,   187,   185,   178,    82,   218,   139,     3,   255,    63,   190,    36,   231,   207,   229,    47,   183,   235,    87,   113,    55,    79,   247,   118,   182,   184,   172,   140,     0,   147,   126,   252,    25,   246,    16,    68,   234,   143,    87,    40,     4,    65,   243,   126,   144,    91,   175,     0,    88,    71,     0,   186,   213,   170,   162,    78,    47,     0,   152,   173,   109,    31,   101,     0,   115,    95,   192,    58,    21,    79,     0,    61,     0,    26,   238,    83,    90,   178,   187,     0,     4,    26,   207,    82,    67,     0,   111,    29,   206,   127,    66,   195,     0),
   (  162,   193,   150,   159,    23,   112,   228,   252,   189,   189,    96,   185,    46,     0,   190,   147,   146,     0,   179,    63,   196,    70,   159,   226,    72,    29,     0,     0,     0,   244,   225,   250,   243,   211,     0,     8,   163,    19,   121,    57,    58,   230,   118,   207,   226,    19,    33,   100,   108,    86,    94,    49,   169,     0,    23,   148,   234,   114,    34,    28,   202,     0,   140,   210,    74,    90,   172,   125,   234,   142,    13,   139,   230,    87,    33,   183,   164,    64,   176,   212,    36,   162,    52,   229,   227,   186,     0,   146,    90,    92,   223,     0,    65,    87,     0,     2,    76,   171,   148,    89,   115,   183,    74,     7,     0,    84,    14,     0,   171,    85,    91,   193,   216,     2,    48,   218,    18,   149,    53,    80,   236,   121,   151,    85,   185,    72,   218,    55),
   (  111,   118,   131,    77,   232,   246,   161,     0,   224,   176,     5,   227,   177,    88,   167,    24,   138,   202,     0,   218,   103,   224,    57,    46,   149,   209,   102,   142,   192,   202,   113,   151,   198,    73,   147,     0,   247,    27,   152,   134,     1,   156,   148,    15,    24,   244,   102,   164,   201,   138,    51,    84,    23,   200,   206,   238,   100,     0,   253,   166,   227,     0,   122,    26,   226,   201,    79,     0,   247,     0,    42,   189,     0,    48,   241,   123,    57,   235,   114,   131,    46,   131,    37,   177,   211,   213,   146,     0,    51,   217,   162,   211,     0,     8,     0,     0,   219,   147,   164,    13,   167,   139,   164,   137,   181,   123,   204,   181,   152,    91,     1,   159,   155,   208,    19,    83,   242,    34,   208,     0,     0,   253,   125,   134,   185,   154,   148,   235),
   (   15,    51,   114,   179,   215,   127,     0,     0,   208,    11,   154,   146,    27,    72,    19,   171,   133,   111,   105,   180,   245,   189,   245,   143,   243,   120,    29,   235,    12,   101,   199,   139,   195,     0,   173,   109,   148,    81,    38,   253,     0,   125,    53,   237,     3,   174,    57,     0,    85,    32,    69,   164,    58,   211,    45,   103,    46,    46,    19,   245,   228,   145,    55,   220,   237,   131,    71,   188,   117,   211,   235,   253,   210,    17,   233,   232,    69,   211,    71,   107,    80,   253,    82,   200,    97,   170,    90,    51,     0,   198,     0,   238,    88,    27,    84,   108,    21,   107,    52,     5,   179,    26,   224,    42,    36,    17,   164,    82,   209,    42,   203,    11,    26,   132,   214,   198,   120,   210,   222,    35,   173,    23,    44,   225,    84,   197,    46,   210),
   (   39,   235,   206,     0,     6,   105,   235,   159,   112,   127,    64,    65,   181,     0,   188,    56,    12,   179,    24,    13,    87,   248,   190,   174,   111,    95,   238,   170,    53,   215,   126,   204,    88,   191,   211,   183,   166,     0,   110,    32,     0,   195,   199,   202,   109,   217,    67,   236,   133,   239,    52,   142,   244,    31,   237,    64,   188,    70,    77,    77,     7,   106,   127,   125,   153,   239,   145,   231,   191,    61,    23,   101,    17,   162,     0,    17,   122,    72,   190,   141,     0,    90,   244,    32,   154,   162,    92,   217,   198,     0,    28,   236,   145,    54,   149,    90,    64,   202,   250,    26,   201,    32,     0,   234,   131,     0,    88,    17,     0,    53,     7,   209,   255,     0,   117,    62,   126,    40,     0,    75,    10,   251,   167,    69,    88,   244,   214,   191),
   (  242,    70,     0,   155,   180,   139,    16,     0,    86,    13,    51,    75,   115,   208,   177,   236,   211,   132,   229,   248,   214,   232,   109,    99,   155,   207,   197,   195,   157,   186,   170,   241,    45,   249,   211,    70,   200,   251,   252,   231,   207,   239,   145,   205,   207,    97,     0,   196,   229,    68,   104,   145,    67,    33,   158,    34,    23,   254,   221,    80,    74,    66,   239,   120,   191,   238,    64,   248,   158,     7,   151,    34,   226,     0,    91,     0,    58,   148,    62,    72,   254,   233,   187,    70,     0,    78,   223,   162,     0,    28,     0,    20,     0,    35,     3,    16,    38,   158,    43,   230,   220,   167,   152,    27,    95,    82,   228,     0,    77,    60,   116,   249,    43,     0,    83,    60,    43,     0,   221,   177,    94,    47,   247,   133,     6,   142,    86,   117),
   (   41,   110,   150,   135,   197,   214,   214,   182,   107,    63,    61,   187,    25,    78,    41,    32,   113,   224,   174,    93,   247,    39,    60,   227,     0,   227,   235,    20,     0,   195,    95,   186,   108,   112,     0,   158,   156,    36,    37,   144,   140,   118,   178,     0,   223,    93,   143,    52,    24,   105,     0,     0,   235,   100,   113,   143,   162,   121,   214,    91,   214,     0,    73,   131,   125,     3,   220,    96,    56,   180,    41,    39,     0,     0,   187,   152,   109,     6,   239,    88,   210,   176,   139,     0,   248,    47,     0,   211,   238,   236,    20,     0,   218,     4,     8,   183,    35,     6,    10,   103,   125,   108,   123,    35,   210,   109,   242,   160,   221,   114,   143,   227,   101,   161,   141,   185,     8,    60,    87,    45,     0,    20,     0,   180,   236,   172,    58,   140),
   (  212,    62,   218,    18,     0,    97,     6,   208,   199,    53,   150,   152,   138,   248,     1,     9,   216,   105,    24,   209,   175,    18,   173,   117,   103,     0,   235,    93,    33,    39,   181,   100,    45,   170,   229,    43,    31,    36,   213,   158,    62,    89,   149,    78,   100,   186,   246,     1,    52,   214,   234,    20,    63,   141,    73,   203,     6,   255,    98,    61,     0,    59,    46,   244,     0,     0,   156,     0,    55,   213,   239,   224,    85,   110,    36,   173,     0,    97,    35,   252,   122,   166,   124,   103,   224,     0,    65,     0,    88,   145,     0,   218,     0,    45,   126,   203,   114,   151,   135,     0,    88,   124,   213,   100,   134,   116,    35,   138,    82,   137,    44,   236,    50,     4,    44,   125,   146,   161,   216,    42,   245,   194,   104,   214,     9,   228,    97,     5),
   (  139,    51,     0,     0,   134,   216,   148,     2,    26,    41,    32,   194,   123,    99,   153,   199,   220,   119,    94,   178,   141,   124,    13,   196,    69,   184,   146,    16,    29,   230,   239,    83,   191,    60,   191,   104,   180,     0,    22,   165,     0,    30,   124,   241,     0,   106,    29,   244,   234,   196,     0,    39,   148,   241,     0,   236,    20,     4,    86,   229,   122,    19,     0,    21,   227,   215,   202,    43,   105,   232,    57,    14,     0,   155,    50,   175,   106,   193,   112,   228,    61,     0,   115,    34,   194,   152,    87,     8,    27,    54,    35,     4,    45,     0,    16,   168,   191,   233,   213,   255,   141,   164,    77,   196,   223,    90,    82,    93,    40,   162,   151,   239,   174,   192,     0,    20,    15,   220,   132,    18,   171,    95,     4,   232,    55,   144,   205,     0),
   (  225,    13,   200,   197,   207,     0,   219,    52,    48,    72,    93,    73,    57,   175,     0,   144,   137,     4,    13,     0,     0,    35,   242,   248,   171,   174,   227,     0,    35,   134,   123,    89,   168,     0,    76,   183,     8,    15,   126,    36,   133,   132,   213,   210,     0,   139,   234,   190,    54,   116,    49,    80,   189,   185,   241,     8,   235,   247,   153,   238,   226,    92,     0,   233,   218,   131,    46,   186,   250,   160,    29,    52,   120,   239,   229,    47,   132,   156,    16,   163,   103,   192,   246,   193,     0,   173,     0,     0,    84,   149,     3,     8,   126,    16,     0,   165,   169,   193,   112,   251,   237,   181,    64,    94,    10,   115,   196,   119,   208,    86,    28,   119,    90,   127,   143,   200,    76,   163,   205,     0,     0,    15,   213,   117,    77,    46,   115,     0),
   (   48,    36,     0,   135,   179,   190,    31,   192,   151,   115,   162,   126,    16,    33,     4,   218,   254,   124,   189,     0,   207,    57,   211,   148,   227,    93,   241,   199,   196,    43,   153,     0,   209,   167,   207,   158,   142,   148,   140,     0,   235,   195,    96,   185,   116,    80,   115,   198,    80,   173,    51,    18,   205,   203,    93,   200,   137,   236,   150,    89,   156,   154,    29,   198,    49,   128,    12,    11,    78,   215,   152,   157,   108,    69,     9,   250,    58,    68,   129,   118,   224,   221,   139,   200,    36,   109,     2,     0,   108,    90,    16,   183,   203,   168,   165,     0,    32,   190,   236,     0,   113,    73,   196,     0,   180,   119,   204,   155,   224,   107,   176,    97,     0,   113,    55,   235,   212,    94,   113,   214,   217,   250,   216,    95,     0,    94,    15,     3),
   (  173,    90,   251,    88,     0,    93,   168,   193,     9,   104,   172,   173,   190,   204,   235,   163,    18,   210,    10,    14,   229,   166,    18,    62,   177,   128,   215,     0,   251,     0,    61,   253,   100,     8,   146,    82,   149,   141,   236,    81,   126,    69,   233,   152,   113,     0,    76,   135,   210,   161,   248,   244,   253,   252,    15,   135,   165,    64,    24,   168,   101,    50,   243,    77,   120,   162,   114,   137,   105,   162,   204,    58,     0,    51,   147,   199,   168,    22,   122,   139,   238,   187,   140,     0,   154,    31,    76,   219,    21,    64,    38,    35,   114,   191,   169,    32,     0,    75,     9,   240,     0,   103,     0,    96,   138,    98,   184,    74,   177,     0,   205,     3,   164,   192,   138,     5,    74,     5,    28,     0,    55,   115,    46,    97,     0,     0,     0,   249),
   (  205,    46,   111,   149,   186,     0,    45,    43,    90,   153,   230,    72,    36,   190,   151,   236,   210,   175,     0,   110,    66,   176,   177,    76,   110,   252,   154,   211,   139,    29,     0,   233,   214,     0,    13,    12,   106,   134,     3,   167,   180,   218,   110,   115,   210,   230,   114,    61,   197,   134,   191,    61,    54,    84,   164,   141,    41,    99,   248,   103,    70,    21,   156,   122,     0,   209,    85,   231,     0,   226,     9,   156,    51,    62,   199,    65,   204,    25,   131,    46,     0,   143,    34,   218,   160,   101,   171,   147,   107,   202,   158,     6,   151,   233,   193,   190,    75,     0,   178,   241,    10,    29,    31,   120,   117,   150,    71,   220,    95,     0,   139,     0,     0,    30,   174,   149,    49,   226,   250,   168,    96,   125,     0,   206,   213,    42,     0,    96),
   (  179,   190,   195,    40,   132,     0,   223,    46,   209,    95,   110,   252,   213,   130,   200,   209,   208,    52,    46,   141,    61,    54,    59,    27,     8,   150,   146,    91,   113,     0,   102,   228,    82,   233,   123,   141,   228,     0,    72,   208,   225,    36,   193,   117,    61,   237,     0,    88,    85,   182,   226,   238,    86,   109,   225,   220,   153,   157,    22,   252,   105,    25,    83,   205,    99,   126,    64,     0,   224,   149,     0,   148,   158,   116,   110,    89,   170,   216,    58,   238,     0,    97,   254,    68,    68,     0,   148,   164,    52,   250,    43,    10,   135,   213,   112,   236,     9,   178,     0,   186,   118,   172,    42,     0,   133,    15,    86,     0,   117,    18,   152,    53,    33,    92,     0,    67,     4,   143,     0,    27,     0,    91,   239,   161,    34,    49,   231,    61),
   (  153,    38,   247,   188,   166,    36,   190,   107,   113,   169,   136,   180,    58,    97,     0,    60,   237,    11,    14,    96,   160,    53,    61,    89,     0,   160,     0,     6,   144,   179,    36,    26,   203,   135,   207,    98,    56,   206,   221,   204,   214,   209,    31,   121,   108,   177,    63,   170,    51,    56,     0,    96,   168,   246,    25,   211,   255,   222,    32,   184,    35,   218,     0,   110,   223,     9,     0,    34,   178,    29,     0,    88,    14,     0,    11,     0,    71,    28,   252,    69,   253,    27,     0,    91,    55,   115,    89,    13,     5,    26,   230,   103,     0,   255,   251,     0,   240,   241,   186,     0,    45,    90,   127,   235,   223,     0,   224,    47,   236,    18,   142,   231,   116,    91,   202,    17,    54,    14,    18,    38,   166,    76,    76,   208,   255,    71,   150,   111),
   (   89,   104,     0,    31,   233,   178,   201,    62,     0,   246,    58,   185,    99,   100,    79,   101,    46,   143,   213,    73,   156,     0,     0,     0,   207,   138,    79,   151,   150,   254,     0,   145,     8,   171,   238,    68,    80,   209,   135,    24,   169,    37,   148,   199,   189,   198,   229,   130,   190,   123,     5,    87,    33,    78,    34,   242,   117,    69,    65,   233,   223,    96,   134,    88,    37,    63,   133,   201,   117,     7,    16,   161,    85,    13,     8,    65,    76,     0,    84,   229,   180,     0,    93,     0,     0,    95,   115,   167,   179,   201,   220,   125,    88,   141,   237,   113,     0,    10,   118,    45,     0,    19,    80,   219,   187,     9,    40,   108,   214,   254,   101,     0,     5,   233,   251,   132,    37,   252,   139,   191,    81,   241,     0,     0,   254,     0,   125,   104),
   (   87,   152,    49,   153,     0,   143,    92,    99,    81,   134,    98,   201,   106,   244,   145,   153,   188,   202,   249,    54,   249,    98,   217,    91,    67,    32,   100,    59,   254,   190,   239,    61,     0,   101,   227,   154,     0,   192,   198,   118,   220,   203,    29,   106,    74,   212,   254,     0,   168,   195,   161,   164,   211,    37,     0,   228,    46,   153,    54,   115,     0,   230,     0,   196,    45,   224,   127,     5,   248,   202,    98,     2,   232,    87,   100,   203,     7,    60,   181,   158,   248,   236,     0,    92,   114,   192,   183,   139,    26,    32,   167,   108,   124,   164,   181,    73,   103,    29,   172,    90,    19,     0,    30,    50,     0,   123,    80,   105,   227,   224,     0,    90,     2,   230,   198,   117,     9,    30,    87,   217,   146,   217,    66,   139,   114,   142,     0,    39),
   (   49,   100,   209,    72,   223,    25,   134,    50,   135,    52,     0,   132,    65,    43,    29,    75,   136,    87,    39,   150,     3,   180,   114,   249,   227,    20,     0,   131,    16,     0,   158,    33,   108,    93,   222,     0,    34,   141,    33,   228,     0,   255,    78,    68,   221,   121,   222,   116,     0,     0,    32,     0,   223,   242,    18,     0,    53,   219,    76,    12,    15,   235,    67,   112,    55,    58,   203,   146,   199,    81,    96,     0,     0,     0,   197,   120,   155,   176,   198,   186,   159,    48,   121,   240,   173,    58,    74,   164,   224,     0,   152,   123,   213,    77,    64,   196,     0,    31,    42,   127,    80,    30,     0,   168,   131,    17,   201,   187,   100,     0,   131,   101,   207,   187,   156,     0,   134,    72,   222,   212,     2,   235,    38,   100,   221,     0,   238,   184),
   (    0,   248,   140,   131,   244,   116,   245,   174,   108,   159,   242,    39,   153,   107,   186,    86,     0,    99,     0,   173,   130,   245,    35,    27,   165,   240,   217,   240,   146,   238,    22,   180,   116,   139,   129,   232,     9,   237,   115,   127,   101,    50,   185,   149,   124,   206,    78,   233,   116,     0,   177,    71,   144,   202,   218,   206,   220,     0,   205,   254,   241,   117,    73,    18,    88,     5,    62,    33,   208,   140,   187,    56,   119,   194,     0,    12,     0,   249,   159,   157,   154,   238,     0,     0,   171,    21,     7,   137,    42,   234,    27,    35,   100,   196,    94,     0,    96,   120,     0,   235,   219,    50,   168,     0,     0,   169,    93,    79,     7,   109,    92,    93,   141,    23,    12,   165,    63,    52,   211,   183,    27,   185,    21,   104,    39,    93,    75,     0),
   (  181,   143,   189,   131,     0,   226,    33,    19,    86,    88,    70,   207,   209,    93,   231,   151,   233,    47,    24,   242,   187,     5,   223,   195,    21,   193,    98,    34,    82,    84,   160,   228,   160,   121,    80,    42,     4,   247,   122,     0,   195,     0,    37,    46,    74,   109,    96,    50,    25,   163,   110,   194,     0,     0,    59,   210,   104,     0,   242,   124,    40,    23,   228,     0,   152,   210,   254,   172,   102,   133,     0,   245,    48,   175,   146,     8,    52,    29,    13,   191,    14,    64,     7,   177,   190,    79,     0,   181,    36,   131,    95,   210,   134,   223,    10,   180,   138,   117,   133,   223,   187,     0,   131,     0,     0,    37,   232,   154,    93,   252,   202,     0,     0,    30,   150,   143,   167,    74,   208,     0,     0,   181,     0,     0,   197,   164,   200,    35),
   (  208,   236,   156,     0,    83,   136,   238,   216,     0,     0,    94,   221,   196,   171,   164,   202,    38,   184,   197,    95,   245,    18,   159,    59,    58,   237,   148,   211,   183,   232,   116,   167,    87,   159,    61,   141,    84,   131,   234,   131,    18,   128,   219,   113,   199,    14,   245,   196,    46,    33,   124,    19,     0,   128,    23,   155,   234,   137,   102,    10,   201,   190,    55,   115,     0,     0,   134,     6,   236,     0,     0,   118,   207,   191,   246,    76,   129,   130,   187,    73,    95,   227,   134,    79,   206,     0,    84,   123,    17,     0,    82,   109,   116,    90,   115,   119,    98,   150,    15,     0,     9,   123,    17,   169,    37,     0,   190,   102,   145,   162,   208,   124,   149,    95,    91,   150,   254,     8,   199,   103,    86,   241,   104,     0,   139,    94,   206,   220),
   (  137,   243,    88,   247,   199,   206,   225,   164,   233,    31,     7,   175,   146,   109,   247,   172,    72,   141,     8,    44,    84,   154,    66,    61,    54,     0,   100,   223,    77,     0,   249,   146,   127,   129,     7,     0,    98,   109,   255,   123,    56,   176,   105,    14,    46,   250,   236,   120,   160,   224,   205,    62,   217,   187,   253,   139,   141,   181,    94,    20,   234,   178,    57,   195,   180,   249,   158,    21,   158,   168,   185,   197,    21,   253,   151,    55,     0,    27,   163,   251,   180,   100,    88,   175,    45,    61,    14,   204,   164,    88,   228,   242,    35,    82,   196,   204,   184,    71,    86,   224,    40,    80,   201,    93,   232,   190,     0,   186,     0,    99,   156,    25,   161,   123,   202,   151,   214,   204,   187,    10,    87,    42,   104,     1,   228,     0,    27,   202),
   (  157,   137,    51,    43,   228,   229,   188,   117,    54,   188,     0,   255,   253,   156,   151,   126,    39,   170,   189,    64,   130,   169,   228,   235,   166,   251,    42,     8,   252,    71,   217,     0,   125,   104,   210,   234,   211,   250,   238,   175,     0,   211,   178,   248,    67,     0,     0,    32,   223,   182,   162,   173,    73,   138,   194,   145,   111,   106,   250,   189,     0,   107,    95,    63,   161,    69,    27,    65,   125,    63,    58,    48,    35,   106,    55,   100,    10,   236,    94,    12,   140,   122,    19,   196,   129,     0,     0,   181,    82,    17,     0,   160,   138,    93,   119,   155,    74,   220,     0,    47,   108,   105,   187,    79,   154,   102,   186,     0,   192,   249,    58,   207,   197,   188,    90,   213,   227,   193,   187,   199,   168,    34,    67,   200,   124,   117,    14,    86),
   (   92,    71,   132,   114,   125,   227,   186,   118,     0,     0,    93,     0,   147,   193,    19,     8,    83,    22,   103,   112,    20,   166,     0,   236,    31,   254,     0,   164,    81,   239,   214,   188,    91,   204,    51,    75,    46,    65,   148,    53,    43,   192,   169,    55,    83,    44,    49,   178,     0,   125,   177,    10,   141,     0,    97,   103,    12,    49,   237,   230,   220,    43,    99,   174,    64,     6,   204,   132,     4,   203,   247,    52,    82,   169,   180,   243,     0,   102,   187,    17,   131,   187,   106,     0,     0,    26,   171,   152,   209,     0,    77,   221,    82,    40,   208,   224,   177,    95,   117,   236,   214,   227,   100,     7,    93,   145,     0,   192,     0,   202,   148,   222,   202,   149,   129,    14,    80,   207,    33,    49,     4,    87,     0,   212,     0,   133,   178,   205),
   (  234,   191,     0,   218,   194,   229,   189,   219,    29,   214,   197,    52,   168,   137,   159,    57,   202,    87,   234,     0,   208,   202,    29,    31,    16,   177,     0,   114,    74,   203,   254,    84,   172,    31,    32,    68,    81,   224,   103,     0,   171,    39,   234,     0,     0,    47,   168,    97,    40,    52,    26,   236,     0,    48,     1,    85,   182,   161,     0,    93,   199,   243,   242,   146,    81,    92,   185,     0,     0,   130,   203,   163,   216,   108,   171,   123,    83,   139,   156,    48,   178,   133,    90,   147,   201,   238,    85,    91,    42,    53,    60,   114,   137,   162,    86,   107,     0,     0,    18,    18,   254,   224,     0,   109,   252,   162,    99,   249,   202,     0,    37,     0,    56,     0,   193,    26,     0,     0,   199,   236,   148,   158,   229,   254,   243,   183,   201,   133),
   (    0,    90,   232,    88,   222,    69,     0,     0,    52,    16,     0,   133,    69,    24,    19,   192,    62,   214,   255,   248,    24,     0,   107,     0,    22,     0,   148,   139,   136,   162,   200,    37,   144,     0,    28,    68,   253,   140,   135,   237,   220,    66,     0,     0,   228,   151,    74,   169,   249,   165,   205,    78,    11,     0,   228,   243,     0,   149,    13,   218,   147,    89,   182,   129,   153,   103,   125,    92,    22,   153,   134,   193,   141,     0,    27,   146,   153,   141,    14,   133,    28,     2,   108,     0,   192,    83,    91,     1,   203,     7,   116,   143,    44,   151,    28,   176,   205,   139,   152,   142,   101,     0,   131,    92,   202,   208,   156,    58,   148,    37,     0,   165,   138,   147,    45,    68,     7,     0,   252,   203,    99,    31,   116,    41,    26,   129,     1,   168),
   (  113,   191,    23,    15,   158,    86,     0,    10,   242,   123,   122,   107,     2,     0,    46,    66,    51,   225,   159,    27,   238,    65,    69,   145,    13,     9,    46,   238,     1,   133,   197,   191,   198,   153,   244,     0,   244,   174,     5,   120,   153,     0,   203,    99,    88,     0,   171,    92,   253,   134,    31,    29,     0,    35,   132,   216,   149,   145,   242,   245,   155,     0,   176,   249,    32,    90,    24,    39,    20,   187,   176,   199,   192,   104,    27,   170,    24,    14,    39,     3,   142,    86,   114,   192,   125,    90,   193,   159,    11,   209,   249,   227,   236,   239,   119,    97,     3,     0,    53,   231,     0,    90,   101,    93,     0,   124,    25,   207,   222,     0,   165,     0,     8,   106,     0,     0,    46,    81,    81,   176,     0,     0,   232,    24,   184,   208,   109,    77),
   (    0,   228,    68,   138,    80,    29,   164,   214,   159,   117,    24,    96,   136,   197,    37,    54,   182,    62,     8,     0,   128,    95,    24,   150,   129,   194,   248,    16,    29,    93,   106,    37,   197,   238,     0,    46,    56,    88,   239,   222,    51,   217,   128,   225,   250,    41,   210,     0,    17,   112,    18,   140,   209,    65,   211,   175,   161,   163,    58,    98,   237,   181,    29,   113,     0,   186,   199,   191,    67,    91,   204,   140,   160,   206,   213,   246,   198,    43,   127,    60,   122,    51,    53,   247,    70,   178,   216,   155,    26,   255,    43,   101,    50,   174,    90,     0,   164,     0,    33,   116,     5,     2,   207,   141,     0,   149,   161,   197,   202,    56,   138,     8,     0,   117,   220,    10,    59,   107,     8,     0,   170,   113,   186,   217,    16,   124,    30,   178),
   (  113,   174,   194,   160,    68,   111,    32,    26,   139,    33,   168,   130,   161,     2,    97,    34,     0,    69,   185,    46,    47,   147,   119,   158,    33,   205,   231,   187,   105,    25,    93,     2,     0,   211,   164,   173,     1,   120,   174,   113,   200,   223,    53,    47,   201,     4,   167,   132,    11,   197,    68,    49,   210,   240,    38,   113,    73,   179,   215,   115,    39,   105,   214,   101,   125,    76,   181,   250,    92,    81,   244,    23,   147,   248,     0,   246,     0,   234,    99,   149,    53,    68,   201,     0,     0,   187,     2,   208,   132,     0,     0,   161,     4,   192,   127,   113,   192,    30,    92,    91,   233,   230,   187,    23,    30,    95,   123,   188,   149,     0,   147,   106,   117,     0,   206,    97,   225,   142,    70,   220,    28,    50,   126,   180,    68,   141,   127,   193),
   (   56,    83,   252,   145,    76,   133,    34,    21,    17,    88,   156,   111,   254,   252,    19,   227,    15,    83,     0,   254,    42,     3,   225,    44,    27,   255,   111,   203,    77,   217,    78,   249,    17,    41,   104,   237,   203,   214,    65,    27,    43,   238,   147,   156,     6,   127,    51,    44,    33,   137,    76,   159,   154,   205,   215,    46,   163,    21,     0,    33,   125,    30,     2,   163,     0,   237,   255,    50,    69,     7,   110,    36,    69,    87,   246,   208,   113,   191,    39,    86,    12,    37,   168,   255,   103,     0,    48,    19,   214,   117,    83,   141,    44,     0,   143,    55,   138,   174,     0,   202,   251,   198,   156,    12,   150,    91,   202,    90,   129,   193,    45,     0,   220,   206,     0,   214,   136,    50,   230,     0,     2,    78,    88,   127,   199,   183,   187,    95),
   (  170,   163,    56,   125,     0,   167,   125,    81,   217,   244,    94,   178,   141,    25,    91,     0,   234,   211,    35,   103,    87,   112,   184,   148,   139,   178,     0,    71,     0,    62,     0,    67,   140,   175,    96,   236,   100,    75,    76,   164,   115,    27,    28,   127,   109,   168,    27,   152,   253,     2,    11,    49,   149,   106,    69,    19,    30,   203,    26,    24,   232,     0,     0,   196,    63,   208,    98,   133,   207,   209,   177,    15,    35,     0,    20,   103,   219,   192,    86,    63,    21,     0,   224,    27,    85,     4,   218,    83,   198,    62,    60,   185,   125,    20,   200,   235,     5,   149,    67,    17,   132,   117,     0,   165,   143,   150,   151,   213,    14,    26,    68,     0,    10,    97,   214,     0,   112,   150,     0,   168,   175,   247,   215,    42,   241,   126,    44,    59),
   (  248,    45,   193,   143,   237,    86,     0,    66,    24,   121,   248,   187,   161,    47,   214,   243,   179,    27,   136,     5,     0,   218,   111,    74,    33,   212,   135,     0,   192,    70,   196,    61,    25,     0,    64,   251,    32,   145,    74,   226,    93,   180,     0,   239,   242,    84,   220,   184,   199,   112,    11,   131,   183,     1,     0,    38,   140,     0,   210,    79,    83,   230,   200,    55,   219,    94,   214,    82,   241,     0,    88,    36,   186,    49,    17,   152,    83,   175,   121,   118,   161,     0,   126,   238,   145,    26,    18,   242,   120,   126,    43,     8,   146,    15,    76,   212,    74,    49,     4,    54,    37,     9,   134,    63,   167,   254,   214,   227,    80,     0,     7,    46,    59,   225,   136,   112,     0,    69,   143,    52,    31,   184,   203,    74,    48,     1,    69,   211),
   (  249,     1,   122,    41,    61,   122,   183,    91,   110,   167,   137,    99,    27,   187,   199,    65,   217,   167,    40,    47,   105,   222,   101,     0,   132,    41,   214,   210,   115,     7,   144,   224,   249,   230,   205,     0,     0,   139,   130,    91,    80,    76,   150,   112,   141,     0,   138,   236,    96,   211,   144,    71,   166,    83,    14,   245,   230,   226,   181,   236,   182,    78,   143,    61,   132,   170,   223,   117,   194,     0,    14,   144,   179,   126,   228,     0,     2,    36,   198,     0,   254,    85,     0,   110,   168,   207,   149,    34,   210,    40,     0,    60,   161,   220,   163,    94,     5,   226,   143,    14,   252,    30,    72,    52,    74,     8,   204,   193,   207,     0,     0,    81,   107,   142,    50,   150,    69,     0,   214,   112,   172,   132,   210,   157,   167,   239,    79,    21),
   (   47,     2,     0,   246,   196,    74,   191,    95,    36,    27,   190,   122,   224,   128,   130,    85,   252,    75,    32,   102,   104,     0,   121,   136,    22,   231,     0,   124,   104,    53,     0,   103,   211,   113,    86,     0,     0,   143,    45,    98,    35,   193,     2,    19,   139,    60,   132,    40,   109,    29,    66,   150,    41,     7,   188,     0,     0,   146,    18,   152,   251,    48,   140,   146,   170,   107,    34,   111,    79,   204,   126,   174,   160,   209,   215,   116,   210,   253,    12,    90,   242,    13,   135,   195,    92,    82,    53,   208,   222,     0,   221,    87,   216,   132,   205,   113,    28,   250,     0,    18,   139,    87,   222,   211,   208,   199,   187,   187,    33,   199,   252,    81,     8,    70,   230,     0,   143,   214,     0,   142,   130,   115,   162,   209,   137,   125,    16,    27),
   (  210,   166,    54,    76,   215,   122,    45,    67,   167,    24,   116,    50,     0,    54,    14,   232,   145,    86,    70,   109,   236,   160,   111,    73,   215,   163,    38,   195,   191,     0,    70,   100,    64,   106,     0,    81,   219,     0,   157,    71,    60,     0,   155,   231,   103,    79,    24,   167,     2,    12,   130,   124,   230,    61,   107,   111,    30,   154,     0,   140,   227,   222,   120,     1,   130,    82,   203,    44,    38,     0,    55,     0,    85,   252,   161,    83,   131,   227,    27,   245,     0,     0,   100,   239,   124,    67,    80,     0,    35,    75,   177,    45,    42,    18,     0,   214,     0,   168,    27,    38,   191,   217,   212,   183,     0,   103,    10,   199,    49,   236,   203,   176,     0,   220,     0,   168,    52,   112,   142,     0,     0,   246,    71,   137,   201,    76,   161,    38),
   (  114,    35,   169,   113,   111,   206,   182,   202,   126,    46,   146,    43,   219,   147,    20,   235,   131,   108,    18,   137,     0,     8,   175,   200,   107,     0,   113,   239,   225,   162,   139,   102,   191,    60,    20,   131,   110,    95,    62,   181,     0,     2,   197,    69,   237,   197,     0,    72,   175,    59,    77,   239,   222,    13,    94,    89,   253,    29,   219,    40,   247,   208,    17,     0,    11,    52,   177,   211,   163,   241,   193,    34,   112,    69,   174,    96,    48,    56,     0,     0,   117,   157,     0,   128,    82,     0,   236,     0,   173,    10,    94,     0,   245,   171,     0,   217,    55,    96,     0,   166,    81,   146,     2,    27,     0,    86,    87,   168,     4,   148,    99,     0,   170,    28,     2,   175,    31,   172,   130,     0,     0,    79,    52,   137,   234,    81,   125,   252),
   (   46,   250,    62,   152,   148,    53,    40,     0,   138,    16,    97,   216,     0,   103,   156,   108,   175,    70,   211,   157,    55,   145,   169,   142,     0,   211,   233,   240,     0,     3,    77,   119,   208,   201,     0,   238,   154,   248,    29,    24,   159,   149,   134,    88,   235,   230,   112,   145,    13,   244,   165,   223,     9,    19,    94,   180,   153,   154,   194,     0,   164,   154,   178,   120,   101,    18,    38,    13,   228,    84,   171,   123,   192,   177,     0,   102,   196,   158,    29,    12,    61,    63,    55,    31,     0,   111,   121,   253,    23,   251,    47,    20,   194,    95,    15,   250,   115,   125,    91,    76,   241,   217,   235,   185,   181,   241,    42,    34,    87,   158,    31,     0,   113,    50,    78,   247,   184,   132,   115,   246,    79,     0,    22,    65,     5,   165,   120,    19),
   (  127,    99,   218,    43,    44,   190,    79,   127,    72,   132,   120,    20,   213,   100,    11,     0,    44,   151,   242,    45,    95,    85,     0,   137,     5,   125,     0,    97,    20,    55,     9,   115,   197,   104,    74,   231,   167,   168,    74,   137,   167,   130,   176,   152,     0,   156,   151,    37,     0,   200,   225,    29,   199,   133,    26,    59,   208,    96,     0,    93,   135,    92,   240,    99,   223,   254,   212,     0,   251,    12,    49,   183,   122,     7,    66,   104,     0,   190,    40,   145,   119,     9,    38,   247,   108,    29,   151,   125,    44,   167,   247,     0,   104,     4,   213,   216,    46,     0,   239,    76,     0,    66,    38,    21,     0,   104,   104,    67,     0,   229,   116,   232,   186,   126,    88,   215,   203,   210,   162,    71,    52,    22,     0,   180,    18,     0,   212,   166),
   (  207,   137,   172,   160,    73,   146,   141,   141,   232,    19,     0,   229,   103,   165,   186,   206,     1,     0,   165,   195,    69,    36,   132,    83,    85,   159,     0,    14,   243,    74,   136,    43,    28,   155,   139,   193,   248,    19,    86,    89,   107,   141,    48,    46,    94,   210,   218,   134,     5,   215,    22,    30,   193,   222,   110,   218,   216,   105,    47,    72,     0,    44,   158,   242,   133,   148,   115,     0,     0,   108,     0,    29,   248,    38,   233,     0,   217,   198,     0,   138,    34,    16,     0,   145,    39,   206,    85,   134,   225,    69,   133,   180,   214,   232,   117,    95,    97,   206,   161,   208,     0,   139,   100,   104,     0,     0,     1,   200,   212,   254,    41,    24,   217,   180,   127,    42,    74,   157,   209,   137,   137,    65,   180,     0,    20,     9,    81,   216),
   (   57,    86,    70,    72,     0,     0,     3,   249,   102,   120,    48,     1,    97,   156,    38,   194,   137,   131,    24,    67,   249,     0,   205,   207,   210,   199,   174,    59,     0,    12,   117,   117,    23,   117,   152,   234,   254,   205,     0,   203,    54,    13,   200,     0,    25,    83,   146,   252,    42,   206,   183,     0,   131,   218,   149,   105,   130,   116,    18,   110,   247,     7,   247,   161,     0,    23,    49,    33,    75,   225,   219,   112,   113,   204,   136,   181,   235,   250,   167,   151,    63,    13,   172,   130,   162,   127,   185,   185,    84,    88,     6,   236,     9,    55,    77,     0,     0,   213,    34,   255,   254,   114,   221,    39,   197,   139,   228,   124,     0,   243,    26,   184,    16,    68,   199,   241,    48,   167,   137,   201,   234,     5,    18,    20,     0,    44,     0,   243),
   (   33,    32,    11,   169,   101,     7,   253,   182,   223,   153,    34,   146,    60,   214,     0,     0,   169,   110,     0,     6,     0,   119,     0,   158,   107,    34,   174,   113,    52,    27,    39,   178,    72,    39,   157,   119,    98,   181,   246,   138,     0,   194,    98,     0,     0,   165,   215,   140,    80,    58,   136,   106,     0,   153,    67,    15,    89,   212,   187,   105,    64,    48,    30,   240,   119,    93,   165,   171,   230,   248,    67,     0,     0,   211,    68,   113,   154,   107,     0,    64,    66,   234,   188,    91,   245,    66,    72,   154,   197,   244,   142,   172,   228,   144,    46,    94,     0,    42,    49,    71,     0,   142,     0,    93,   164,    94,     0,   117,   133,   183,   129,   208,   124,   141,   183,   126,     1,   239,   125,    76,    81,   165,     0,     9,    44,     0,   227,   252),
   (  139,   214,   137,    48,     0,   255,   212,   132,    59,    25,    54,   173,     0,    72,    95,    56,     0,    52,   152,    64,   122,   149,   101,     0,    99,    74,   231,   244,     5,     0,    72,     0,   246,   176,    57,    79,   152,    98,   169,    51,   143,   152,   221,   218,     8,    42,   135,   117,   167,    51,     2,     1,    81,    13,    85,    15,    85,     1,    86,   185,    36,    25,   159,   240,    20,   227,   134,    22,   165,   243,   170,     0,     0,   251,   232,   180,   240,     3,   121,    84,    75,   132,   239,   210,   177,   195,   218,   148,    46,   214,    86,    58,    97,   205,   115,    15,     0,     0,   231,   150,   125,     0,   238,    75,   200,   206,    27,    14,   178,   201,     1,   109,    30,   127,   187,    44,    69,    79,    16,   161,   125,   120,   212,    81,     0,   227,     0,   150),
   (  214,   240,    97,   105,   254,     0,   192,    61,    80,   249,     0,   195,     0,    33,   125,   130,   134,   162,    72,   253,   107,   213,   212,   216,   252,   169,   231,     0,     0,    99,   165,   191,   245,     0,   151,    96,     6,   219,   169,    86,   236,    28,    27,   148,    23,   133,   253,     0,   243,    36,   237,    24,     0,   169,   196,    63,   222,   184,    16,   187,   101,     0,   196,   208,    83,   155,   250,    34,   181,     4,   107,    98,   157,     0,    41,   106,   122,   115,   250,   206,   163,     4,   246,    52,     0,     0,    55,   235,   210,   191,   117,   140,     5,     0,     0,     3,   249,    96,    61,   111,   104,    39,   184,     0,    35,   220,   202,    86,   205,   133,   168,    77,   178,   193,    95,    59,   211,    21,    27,    38,   252,    19,   166,   216,   243,   252,   150,     0));
   
  type key is array(0 to 127) of integer;
  constant answer_key : key :=
  ( 0, 7733260, 458760, 4980753, 5, 851980, 8126477, 5, 5177365, 5767193, 5308432, 1769481, 7274512, 7405577, 6029324, 131087, 8060948, 4456464, 1376271, 3342346, 3670026, 8, 262154, 1, 7995408, 1376274, 3080210, 458758, 8257551, 5505039, 1507338, 7405577, 131082, 3997711, 4587535, 3932174, 7405576, 2686982, 7274515, 131083, 5701645, 2949124, 1769480, 2359306, 4194315, 1507331, 1376266, 6029324, 2097166, 4521997, 8257548, 458761, 262153, 1441808, 7, 262150, 7, 6094859, 1769488, 2293778, 4063244, 131084, 7471114, 458764, 8, 5963790, 3080205, 65551, 7077902, 1769483, 1310731, 2031629, 2097164, 2424843, 6225940, 2424841, 3538958, 8257549, 2949139, 851979, 4521996, 7208973, 2555916, 2686982, 11, 2752523, 7405577, 7208972, 2883598, 262155, 8126480, 6094859, 7405579, 458759, 3604494, 5636107, 7274513, 5963793, 7602195, 1769484, 3276817, 4653071, 7864328, 5636112, 2359308, 2949137, 8060948, 1769486, 7864330, 3538952, 8257547, 5177358, 6619153, 2949127, 7864328, 5570575, 1245199, 65549, 2752522, 4128781, 2686982, 8126479, 6094859, 3145747, 720906, 1245200, 3342346, 2359310 );

  constant TEST_SIZE : integer := 128;
  constant MAX_CYCLES : integer  := TEST_SIZE*4;

  signal clk : std_logic := '0';
  signal rst : std_logic := '1';

  signal mmap_wr_en   : std_logic                         := '0';
  signal mmap_wr_addr : std_logic_vector(MMAP_ADDR_RANGE) := (others => '0');
  signal mmap_wr_data : std_logic_vector(MMAP_DATA_RANGE) := (others => '0');

  signal mmap_rd_en   : std_logic                         := '0';
  signal mmap_rd_addr : std_logic_vector(MMAP_ADDR_RANGE) := (others => '0');
  signal mmap_rd_data : std_logic_vector(MMAP_DATA_RANGE);

  signal sim_done : std_logic := '0';

begin

  UUT : entity work.user_app
    port map (
      clk          => clk,
      rst          => rst,
      mmap_wr_en   => mmap_wr_en,
      mmap_wr_addr => mmap_wr_addr,
      mmap_wr_data => mmap_wr_data,
      mmap_rd_en   => mmap_rd_en,
      mmap_rd_addr => mmap_rd_addr,
      mmap_rd_data => mmap_rd_data);

  -- toggle clock
  clk <= not clk after 5 ns when sim_done = '0' else clk;

  -- process to test different inputs
  process

    procedure clearMMAP is
    begin
      mmap_rd_en <= '0';
      mmap_wr_en <= '0';
    end clearMMAP;

    variable errors : integer := 0;

    variable result : std_logic_vector(C_MMAP_DATA_WIDTH-1 downto 0);
    variable done   : std_logic;
    variable count  : integer;

  begin
    report "============================SIMULATION START============================" severity note;
    -- reset circuit  
    rst <= '1';
    clearMMAP;
    wait for 200 ns;

    rst <= '0';
    wait until clk'event and clk = '1';
    wait until clk'event and clk = '1';

    -- write contents to input ram, which starts at addr 0
    for i in 0 to (TEST_SIZE / 4) - 1 loop
      mmap_wr_addr <= C_MEM_IN_SEL_ADDR;
      mmap_wr_en   <= '1';
      mmap_wr_data <= std_logic_vector(to_unsigned(i, C_MMAP_DATA_WIDTH));
      wait until clk'event and clk = '1';
      clearMMAP;
      for j in 0 to TEST_SIZE - 1 loop
        mmap_wr_addr <= std_logic_vector(to_unsigned(j, C_MMAP_ADDR_WIDTH));
        mmap_wr_en   <= '1';
        mmap_wr_data <= std_logic_vector(to_unsigned(input_key(4*i, j), 8) &
                                         to_unsigned(input_key(4*i+1, j), 8) &
                                         to_unsigned(input_key(4*i+2, j), 8) &
                                         to_unsigned(input_key(4*i+3, j), 8));
        wait until clk'event and clk = '1';
        clearMMAP;
      end loop;      
    end loop;

    -- send size
    mmap_wr_addr <= C_SIZE_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(TEST_SIZE, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;

    -- send src
    mmap_wr_addr <= C_SRC_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(0, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;

    ---- send go = 1 over memory map
    mmap_wr_addr <= C_GO_ADDR;
    mmap_wr_en   <= '1';
    mmap_wr_data <= std_logic_vector(to_unsigned(1, C_MMAP_DATA_WIDTH));
    wait until clk'event and clk = '1';
    clearMMAP;
    
    done  := '0';
    count := 0;

    -- read the done signal every cycle to see if the circuit has
    -- completed.
    --
    -- equivalent to wait until (done = '1') for TIMEOUT;      
    while done = '0' and count < MAX_CYCLES loop

      mmap_rd_addr <= C_DONE_ADDR;
      mmap_rd_en   <= '1';
      wait until clk'event and clk = '1';
      clearMMAP;
      -- give entity one cycle to respond
      wait until clk'event and clk = '1';
      done         := mmap_rd_data(0);
      count        := count + 1;
    end loop;

    if (done /= '1') then
      errors := errors + 1;
      report "Done signal not asserted before timeout.";
    end if;

    -- read outputs from output memory
    for i in 0 to TEST_SIZE-1 loop
      mmap_rd_addr   <= std_logic_vector(to_unsigned(i, C_MMAP_ADDR_WIDTH));
      mmap_rd_en     <= '1';            
      wait until clk'event and clk = '1';
      clearMMAP;
      -- give entity one cycle to respond
      wait until clk'event and clk = '1';
      result := mmap_rd_data;

      if (unsigned(result) /= answer_key(i)) then
        errors := errors + 1;
        report "Result for " & integer'image(i) &
          " is incorrect. The output is " &
          integer'image(to_integer(unsigned(result))) &
          " but should be " & integer'image(answer_key(i));
      end if;
    end loop;  -- i

    report "SIMULATION FINISHED!!!";
    report "TOTAL ERRORS : " & integer'image(errors);
    report "=============================SIMULATION END=============================" severity note;
    sim_done <= '1';
    wait;

  end process;
end tb;
