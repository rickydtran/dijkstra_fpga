../ip_repo/accelerator_1.0/src/comp_lt.vhd